`include "coherence_controller_if.vh"

module coherence_controller(
	coherence_controller_if.cc ccif
);

endmodule
