// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "02/01/2017 17:00:06"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	CLK,
	nRST,
	\syif.halt ,
	\syif.load ,
	\syif.addr ,
	\syif.store ,
	\syif.REN ,
	\syif.WEN ,
	\syif.tbCTRL );
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	CLK;
input 	nRST;
output 	\syif.halt ;
output 	[31:0] \syif.load ;
input 	[31:0] \syif.addr ;
input 	[31:0] \syif.store ;
input 	\syif.REN ;
input 	\syif.WEN ;
input 	\syif.tbCTRL ;

// Design Ports Information
// syif.halt	=>  Location: PIN_T7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[0]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[1]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[2]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[3]	=>  Location: PIN_G22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[4]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[5]	=>  Location: PIN_G19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[6]	=>  Location: PIN_J15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[7]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[8]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[9]	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[10]	=>  Location: PIN_G20,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[11]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[12]	=>  Location: PIN_C16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[13]	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[14]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[15]	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[16]	=>  Location: PIN_R2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[17]	=>  Location: PIN_R6,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[18]	=>  Location: PIN_A10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[19]	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[20]	=>  Location: PIN_AB12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[21]	=>  Location: PIN_A11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[22]	=>  Location: PIN_P2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[23]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[24]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[25]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[26]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[27]	=>  Location: PIN_H21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[28]	=>  Location: PIN_J16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[29]	=>  Location: PIN_N8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[30]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[31]	=>  Location: PIN_A12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// nRST	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.tbCTRL	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[1]	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[0]	=>  Location: PIN_G13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[3]	=>  Location: PIN_M2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[2]	=>  Location: PIN_P1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[5]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[4]	=>  Location: PIN_H13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[7]	=>  Location: PIN_B18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[6]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[9]	=>  Location: PIN_J13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[8]	=>  Location: PIN_E14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[11]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[10]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[13]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[12]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[15]	=>  Location: PIN_R22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[14]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[17]	=>  Location: PIN_R1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[16]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[19]	=>  Location: PIN_M23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[18]	=>  Location: PIN_AB13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[21]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[20]	=>  Location: PIN_D10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[23]	=>  Location: PIN_F17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[22]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[25]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[24]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[27]	=>  Location: PIN_B11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[26]	=>  Location: PIN_B10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[29]	=>  Location: PIN_R23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[28]	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[31]	=>  Location: PIN_J12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[30]	=>  Location: PIN_R7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.WEN	=>  Location: PIN_R21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.REN	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// CLK	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[0]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[1]	=>  Location: PIN_H16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[2]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[3]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[4]	=>  Location: PIN_H19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[5]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[6]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[7]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[8]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[9]	=>  Location: PIN_H17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[10]	=>  Location: PIN_N21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[11]	=>  Location: PIN_AF17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[12]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[13]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[14]	=>  Location: PIN_P21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[15]	=>  Location: PIN_G18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[16]	=>  Location: PIN_G14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[17]	=>  Location: PIN_R3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[18]	=>  Location: PIN_D16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[19]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[20]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[21]	=>  Location: PIN_AC11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[22]	=>  Location: PIN_AB16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[23]	=>  Location: PIN_AE14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[24]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[25]	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[26]	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[27]	=>  Location: PIN_E17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[28]	=>  Location: PIN_G16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[29]	=>  Location: PIN_P25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[30]	=>  Location: PIN_J17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[31]	=>  Location: PIN_P26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tms	=>  Location: PIN_P8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tck	=>  Location: PIN_P5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdi	=>  Location: PIN_P7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdo	=>  Location: PIN_P6,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ;
wire \CPU|DP|dpif.halt~_Duplicate_1_q ;
wire \RAM|ramif.ramload[0]~0_combout ;
wire \RAM|LessThan1~0_combout ;
wire \CPU|DP|ru|ruif.dWEN_r~q ;
wire \CPU|DP|ru|ruif.dREN_r~q ;
wire \ramaddr~0_combout ;
wire \ramaddr~1_combout ;
wire \ramaddr~2_combout ;
wire \ramaddr~3_combout ;
wire \ramaddr~4_combout ;
wire \ramaddr~5_combout ;
wire \ramaddr~6_combout ;
wire \ramaddr~7_combout ;
wire \ramaddr~8_combout ;
wire \ramaddr~9_combout ;
wire \ramaddr~10_combout ;
wire \ramaddr~11_combout ;
wire \ramaddr~12_combout ;
wire \ramaddr~13_combout ;
wire \ramaddr~14_combout ;
wire \ramaddr~15_combout ;
wire \RAM|always0~4_combout ;
wire \ramaddr~16_combout ;
wire \ramaddr~17_combout ;
wire \ramaddr~18_combout ;
wire \ramaddr~19_combout ;
wire \ramaddr~20_combout ;
wire \ramaddr~21_combout ;
wire \ramaddr~22_combout ;
wire \ramaddr~23_combout ;
wire \ramaddr~24_combout ;
wire \ramaddr~25_combout ;
wire \ramaddr~26_combout ;
wire \ramaddr~27_combout ;
wire \ramaddr~28_combout ;
wire \ramaddr~29_combout ;
wire \ramaddr~30_combout ;
wire \ramaddr~31_combout ;
wire \RAM|always0~9_combout ;
wire \ramaddr~32_combout ;
wire \ramaddr~33_combout ;
wire \ramaddr~34_combout ;
wire \ramaddr~35_combout ;
wire \ramaddr~36_combout ;
wire \ramaddr~37_combout ;
wire \ramaddr~38_combout ;
wire \ramaddr~39_combout ;
wire \ramaddr~40_combout ;
wire \ramaddr~41_combout ;
wire \ramaddr~42_combout ;
wire \ramaddr~43_combout ;
wire \ramaddr~44_combout ;
wire \ramaddr~45_combout ;
wire \ramaddr~46_combout ;
wire \ramaddr~47_combout ;
wire \ramaddr~48_combout ;
wire \ramaddr~49_combout ;
wire \ramaddr~50_combout ;
wire \ramaddr~51_combout ;
wire \ramaddr~52_combout ;
wire \ramaddr~53_combout ;
wire \ramaddr~54_combout ;
wire \ramaddr~55_combout ;
wire \ramaddr~56_combout ;
wire \ramaddr~57_combout ;
wire \ramaddr~58_combout ;
wire \ramaddr~59_combout ;
wire \ramaddr~60_combout ;
wire \ramaddr~61_combout ;
wire \ramaddr~62_combout ;
wire \ramaddr~63_combout ;
wire \ramWEN~0_combout ;
wire \ramREN~0_combout ;
wire \ramREN~1_combout ;
wire \RAM|always0~20_combout ;
wire \RAM|always0~21_combout ;
wire \RAM|ramif.ramload[0]~1_combout ;
wire \RAM|always1~1_combout ;
wire \RAM|ramif.ramload[1]~2_combout ;
wire \RAM|ramif.ramload[2]~3_combout ;
wire \RAM|ramif.ramload[2]~4_combout ;
wire \RAM|ramif.ramload[3]~5_combout ;
wire \RAM|ramif.ramload[4]~6_combout ;
wire \RAM|ramif.ramload[4]~7_combout ;
wire \RAM|ramif.ramload[5]~8_combout ;
wire \RAM|ramif.ramload[5]~9_combout ;
wire \RAM|ramif.ramload[6]~10_combout ;
wire \RAM|ramif.ramload[7]~11_combout ;
wire \RAM|ramif.ramload[8]~12_combout ;
wire \RAM|ramif.ramload[9]~13_combout ;
wire \RAM|ramif.ramload[10]~14_combout ;
wire \RAM|ramif.ramload[11]~15_combout ;
wire \RAM|ramif.ramload[12]~16_combout ;
wire \RAM|ramif.ramload[13]~17_combout ;
wire \RAM|ramif.ramload[14]~18_combout ;
wire \RAM|ramif.ramload[15]~19_combout ;
wire \RAM|ramif.ramload[16]~20_combout ;
wire \RAM|ramif.ramload[16]~21_combout ;
wire \RAM|ramif.ramload[17]~22_combout ;
wire \RAM|ramif.ramload[17]~23_combout ;
wire \RAM|ramif.ramload[18]~24_combout ;
wire \RAM|ramif.ramload[19]~25_combout ;
wire \RAM|ramif.ramload[20]~26_combout ;
wire \RAM|ramif.ramload[21]~27_combout ;
wire \RAM|ramif.ramload[22]~28_combout ;
wire \RAM|ramif.ramload[23]~29_combout ;
wire \RAM|ramif.ramload[24]~30_combout ;
wire \RAM|ramif.ramload[25]~31_combout ;
wire \RAM|ramif.ramload[26]~32_combout ;
wire \RAM|ramif.ramload[26]~33_combout ;
wire \RAM|ramif.ramload[27]~34_combout ;
wire \RAM|ramif.ramload[27]~35_combout ;
wire \RAM|ramif.ramload[28]~36_combout ;
wire \RAM|ramif.ramload[28]~37_combout ;
wire \RAM|ramif.ramload[29]~38_combout ;
wire \RAM|ramif.ramload[29]~39_combout ;
wire \RAM|ramif.ramload[30]~40_combout ;
wire \RAM|ramif.ramload[30]~41_combout ;
wire \RAM|ramif.ramload[31]~42_combout ;
wire \RAM|ramif.ramload[31]~43_combout ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ;
wire \CPUCLK~q ;
wire \CPU|DP|rf|Mux63~9_combout ;
wire \CPU|DP|rf|Mux63~19_combout ;
wire \CPU|CM|dcif.imemload[20]~10_combout ;
wire \ramstore~0_combout ;
wire \ramstore~1_combout ;
wire \CPU|DP|rf|Mux33~9_combout ;
wire \CPU|DP|rf|Mux33~19_combout ;
wire \CPU|DP|rf|Mux34~9_combout ;
wire \CPU|DP|rf|Mux34~19_combout ;
wire \CPU|DP|rf|Mux35~9_combout ;
wire \CPU|DP|rf|Mux35~19_combout ;
wire \CPU|DP|rf|Mux36~9_combout ;
wire \CPU|DP|rf|Mux36~19_combout ;
wire \CPU|DP|rf|Mux37~9_combout ;
wire \CPU|DP|rf|Mux37~19_combout ;
wire \CPU|DP|rf|Mux38~9_combout ;
wire \CPU|DP|rf|Mux38~19_combout ;
wire \CPU|DP|rf|Mux39~9_combout ;
wire \CPU|DP|rf|Mux39~19_combout ;
wire \CPU|DP|rf|Mux40~9_combout ;
wire \CPU|DP|rf|Mux40~19_combout ;
wire \CPU|DP|rf|Mux41~9_combout ;
wire \CPU|DP|rf|Mux41~19_combout ;
wire \CPU|DP|rf|Mux42~9_combout ;
wire \CPU|DP|rf|Mux42~19_combout ;
wire \CPU|DP|rf|Mux43~9_combout ;
wire \CPU|DP|rf|Mux43~19_combout ;
wire \CPU|DP|rf|Mux44~9_combout ;
wire \CPU|DP|rf|Mux44~19_combout ;
wire \CPU|DP|rf|Mux45~9_combout ;
wire \CPU|DP|rf|Mux45~19_combout ;
wire \CPU|DP|rf|Mux46~9_combout ;
wire \CPU|DP|rf|Mux46~19_combout ;
wire \CPU|DP|rf|Mux47~9_combout ;
wire \CPU|DP|rf|Mux47~19_combout ;
wire \CPU|DP|rf|Mux48~9_combout ;
wire \CPU|DP|rf|Mux48~19_combout ;
wire \CPU|DP|rf|Mux49~9_combout ;
wire \CPU|DP|rf|Mux49~19_combout ;
wire \CPU|DP|rf|Mux50~9_combout ;
wire \CPU|DP|rf|Mux50~19_combout ;
wire \CPU|DP|rf|Mux51~9_combout ;
wire \CPU|DP|rf|Mux51~19_combout ;
wire \CPU|DP|rf|Mux52~9_combout ;
wire \CPU|DP|rf|Mux52~19_combout ;
wire \CPU|DP|rf|Mux53~9_combout ;
wire \CPU|DP|rf|Mux53~19_combout ;
wire \CPU|DP|rf|Mux54~9_combout ;
wire \CPU|DP|rf|Mux54~19_combout ;
wire \CPU|DP|rf|Mux55~9_combout ;
wire \CPU|DP|rf|Mux55~19_combout ;
wire \CPU|DP|rf|Mux56~9_combout ;
wire \CPU|DP|rf|Mux56~19_combout ;
wire \CPU|DP|rf|Mux57~9_combout ;
wire \CPU|DP|rf|Mux57~19_combout ;
wire \CPU|DP|rf|Mux58~9_combout ;
wire \CPU|DP|rf|Mux58~19_combout ;
wire \CPU|DP|rf|Mux59~9_combout ;
wire \CPU|DP|rf|Mux59~19_combout ;
wire \CPU|DP|rf|Mux60~9_combout ;
wire \CPU|DP|rf|Mux60~19_combout ;
wire \CPU|DP|rf|Mux61~9_combout ;
wire \CPU|DP|rf|Mux61~19_combout ;
wire \CPU|DP|rf|Mux62~9_combout ;
wire \CPU|DP|rf|Mux62~19_combout ;
wire \CPU|DP|rf|Mux32~9_combout ;
wire \CPU|DP|rf|Mux32~19_combout ;
wire \ramstore~2_combout ;
wire \ramstore~3_combout ;
wire \ramstore~4_combout ;
wire \ramstore~5_combout ;
wire \ramstore~6_combout ;
wire \ramstore~7_combout ;
wire \ramstore~8_combout ;
wire \ramstore~9_combout ;
wire \ramstore~10_combout ;
wire \ramstore~11_combout ;
wire \ramstore~12_combout ;
wire \ramstore~13_combout ;
wire \ramstore~14_combout ;
wire \ramstore~15_combout ;
wire \ramstore~16_combout ;
wire \ramstore~17_combout ;
wire \ramstore~18_combout ;
wire \ramstore~19_combout ;
wire \ramstore~20_combout ;
wire \ramstore~21_combout ;
wire \ramstore~22_combout ;
wire \ramstore~23_combout ;
wire \ramstore~24_combout ;
wire \ramstore~25_combout ;
wire \ramstore~26_combout ;
wire \ramstore~27_combout ;
wire \ramstore~28_combout ;
wire \ramstore~29_combout ;
wire \ramstore~30_combout ;
wire \ramstore~31_combout ;
wire \ramstore~32_combout ;
wire \ramstore~33_combout ;
wire \ramstore~34_combout ;
wire \ramstore~35_combout ;
wire \ramstore~36_combout ;
wire \ramstore~37_combout ;
wire \ramstore~38_combout ;
wire \ramstore~39_combout ;
wire \ramstore~40_combout ;
wire \ramstore~41_combout ;
wire \ramstore~42_combout ;
wire \ramstore~43_combout ;
wire \ramstore~44_combout ;
wire \ramstore~45_combout ;
wire \ramstore~46_combout ;
wire \ramstore~47_combout ;
wire \ramstore~48_combout ;
wire \ramstore~49_combout ;
wire \ramstore~50_combout ;
wire \ramstore~51_combout ;
wire \ramstore~52_combout ;
wire \ramstore~53_combout ;
wire \ramstore~54_combout ;
wire \ramstore~55_combout ;
wire \ramstore~56_combout ;
wire \ramstore~57_combout ;
wire \ramstore~58_combout ;
wire \ramstore~59_combout ;
wire \ramstore~60_combout ;
wire \ramstore~61_combout ;
wire \ramstore~62_combout ;
wire \ramstore~63_combout ;
wire \Equal0~0_combout ;
wire \CPUCLK~0_combout ;
wire \count[3]~0_combout ;
wire \count[2]~1_combout ;
wire \count[1]~2_combout ;
wire \count~3_combout ;
wire \ramaddr~29_wirecell_combout ;
wire \altera_internal_jtag~TCKUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~10 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
wire \nRST~input_o ;
wire \syif.tbCTRL~input_o ;
wire \syif.addr[1]~input_o ;
wire \syif.addr[0]~input_o ;
wire \syif.addr[3]~input_o ;
wire \syif.addr[2]~input_o ;
wire \syif.addr[5]~input_o ;
wire \syif.addr[4]~input_o ;
wire \syif.addr[7]~input_o ;
wire \syif.addr[6]~input_o ;
wire \syif.addr[9]~input_o ;
wire \syif.addr[8]~input_o ;
wire \syif.addr[11]~input_o ;
wire \syif.addr[10]~input_o ;
wire \syif.addr[13]~input_o ;
wire \syif.addr[12]~input_o ;
wire \syif.addr[15]~input_o ;
wire \syif.addr[14]~input_o ;
wire \syif.addr[17]~input_o ;
wire \syif.addr[16]~input_o ;
wire \syif.addr[19]~input_o ;
wire \syif.addr[18]~input_o ;
wire \syif.addr[21]~input_o ;
wire \syif.addr[20]~input_o ;
wire \syif.addr[23]~input_o ;
wire \syif.addr[22]~input_o ;
wire \syif.addr[25]~input_o ;
wire \syif.addr[24]~input_o ;
wire \syif.addr[27]~input_o ;
wire \syif.addr[26]~input_o ;
wire \syif.addr[29]~input_o ;
wire \syif.addr[28]~input_o ;
wire \syif.addr[31]~input_o ;
wire \syif.addr[30]~input_o ;
wire \syif.WEN~input_o ;
wire \syif.REN~input_o ;
wire \CLK~input_o ;
wire \syif.store[0]~input_o ;
wire \syif.store[1]~input_o ;
wire \syif.store[2]~input_o ;
wire \syif.store[3]~input_o ;
wire \syif.store[4]~input_o ;
wire \syif.store[5]~input_o ;
wire \syif.store[6]~input_o ;
wire \syif.store[7]~input_o ;
wire \syif.store[8]~input_o ;
wire \syif.store[9]~input_o ;
wire \syif.store[10]~input_o ;
wire \syif.store[11]~input_o ;
wire \syif.store[12]~input_o ;
wire \syif.store[13]~input_o ;
wire \syif.store[14]~input_o ;
wire \syif.store[15]~input_o ;
wire \syif.store[16]~input_o ;
wire \syif.store[17]~input_o ;
wire \syif.store[18]~input_o ;
wire \syif.store[19]~input_o ;
wire \syif.store[20]~input_o ;
wire \syif.store[21]~input_o ;
wire \syif.store[22]~input_o ;
wire \syif.store[23]~input_o ;
wire \syif.store[24]~input_o ;
wire \syif.store[25]~input_o ;
wire \syif.store[26]~input_o ;
wire \syif.store[27]~input_o ;
wire \syif.store[28]~input_o ;
wire \syif.store[29]~input_o ;
wire \syif.store[30]~input_o ;
wire \syif.store[31]~input_o ;
wire \altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire \CPUCLK~clkctrl_outclk ;
wire \nRST~inputclkctrl_outclk ;
wire \CLK~inputclkctrl_outclk ;
wire \CPU|DP|dpif.halt~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TDIUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
wire [9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
wire [5:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
wire [15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
wire [3:0] count;
wire [31:0] \CPU|DP|PC ;
wire [31:0] \CPU|CM|daddr ;
wire [3:0] \RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg ;


ram RAM(
	.is_in_use_reg(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.LessThan1(\RAM|LessThan1~0_combout ),
	.ramaddr(\ramaddr~1_combout ),
	.ramaddr1(\ramaddr~3_combout ),
	.ramaddr2(\ramaddr~5_combout ),
	.ramaddr3(\ramaddr~7_combout ),
	.ramaddr4(\ramaddr~9_combout ),
	.ramaddr5(\ramaddr~11_combout ),
	.ramaddr6(\ramaddr~13_combout ),
	.ramaddr7(\ramaddr~15_combout ),
	.always0(\RAM|always0~4_combout ),
	.ramaddr8(\ramaddr~17_combout ),
	.ramaddr9(\ramaddr~19_combout ),
	.ramaddr10(\ramaddr~21_combout ),
	.ramaddr11(\ramaddr~23_combout ),
	.ramaddr12(\ramaddr~25_combout ),
	.ramaddr13(\ramaddr~27_combout ),
	.ramaddr14(\ramaddr~29_combout ),
	.ramaddr15(\ramaddr~31_combout ),
	.always01(\RAM|always0~9_combout ),
	.ramaddr16(\ramaddr~33_combout ),
	.ramaddr17(\ramaddr~35_combout ),
	.\ramif.ramaddr ({\ramaddr~61_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\ramaddr~37_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.ramaddr18(\ramaddr~39_combout ),
	.ramaddr19(\ramaddr~41_combout ),
	.ramaddr20(\ramaddr~43_combout ),
	.ramaddr21(\ramaddr~45_combout ),
	.ramaddr22(\ramaddr~47_combout ),
	.ramaddr23(\ramaddr~49_combout ),
	.ramaddr24(\ramaddr~51_combout ),
	.ramaddr25(\ramaddr~53_combout ),
	.ramaddr26(\ramaddr~55_combout ),
	.ramaddr27(\ramaddr~57_combout ),
	.ramaddr28(\ramaddr~59_combout ),
	.ramaddr29(\ramaddr~63_combout ),
	.\ramif.ramWEN (\ramWEN~0_combout ),
	.\ramif.ramREN (\ramREN~1_combout ),
	.always02(\RAM|always0~20_combout ),
	.always03(\RAM|always0~21_combout ),
	.ramiframload_01(\RAM|ramif.ramload[0]~1_combout ),
	.always1(\RAM|always1~1_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~2_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~3_combout ),
	.ramiframload_21(\RAM|ramif.ramload[2]~4_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~5_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~6_combout ),
	.ramiframload_41(\RAM|ramif.ramload[4]~7_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~8_combout ),
	.ramiframload_51(\RAM|ramif.ramload[5]~9_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~10_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~11_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~12_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~13_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~14_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~15_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~16_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~17_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~18_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~19_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~20_combout ),
	.ramiframload_161(\RAM|ramif.ramload[16]~21_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~22_combout ),
	.ramiframload_171(\RAM|ramif.ramload[17]~23_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~24_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~25_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~26_combout ),
	.ramiframload_211(\RAM|ramif.ramload[21]~27_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~28_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~29_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~30_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~31_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~32_combout ),
	.ramiframload_261(\RAM|ramif.ramload[26]~33_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~34_combout ),
	.ramiframload_271(\RAM|ramif.ramload[27]~35_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~36_combout ),
	.ramiframload_281(\RAM|ramif.ramload[28]~37_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~38_combout ),
	.ramiframload_291(\RAM|ramif.ramload[29]~39_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~40_combout ),
	.ramiframload_301(\RAM|ramif.ramload[30]~41_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~42_combout ),
	.ramiframload_311(\RAM|ramif.ramload[31]~43_combout ),
	.ir_loaded_address_reg_0(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.ir_loaded_address_reg_1(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.ir_loaded_address_reg_2(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.ir_loaded_address_reg_3(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.tdo(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.ramstore(\ramstore~1_combout ),
	.ramstore1(\ramstore~3_combout ),
	.ramstore2(\ramstore~5_combout ),
	.ramstore3(\ramstore~7_combout ),
	.ramstore4(\ramstore~9_combout ),
	.ramstore5(\ramstore~11_combout ),
	.ramstore6(\ramstore~13_combout ),
	.ramstore7(\ramstore~15_combout ),
	.ramstore8(\ramstore~17_combout ),
	.ramstore9(\ramstore~19_combout ),
	.ramstore10(\ramstore~21_combout ),
	.ramstore11(\ramstore~23_combout ),
	.ramstore12(\ramstore~25_combout ),
	.ramstore13(\ramstore~27_combout ),
	.ramstore14(\ramstore~29_combout ),
	.ramstore15(\ramstore~31_combout ),
	.ramstore16(\ramstore~33_combout ),
	.ramstore17(\ramstore~35_combout ),
	.ramstore18(\ramstore~37_combout ),
	.ramstore19(\ramstore~39_combout ),
	.ramstore20(\ramstore~41_combout ),
	.ramstore21(\ramstore~43_combout ),
	.ramstore22(\ramstore~45_combout ),
	.ramstore23(\ramstore~47_combout ),
	.ramstore24(\ramstore~49_combout ),
	.ramstore25(\ramstore~51_combout ),
	.ramstore26(\ramstore~53_combout ),
	.ramstore27(\ramstore~55_combout ),
	.ramstore28(\ramstore~57_combout ),
	.ramstore29(\ramstore~59_combout ),
	.ramstore30(\ramstore~61_combout ),
	.ramstore31(\ramstore~63_combout ),
	.ramaddr30(\ramaddr~29_wirecell_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.irf_reg_0_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.node_ena_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.clr_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.virtual_ir_scan_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.state_5(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.state_8(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.nRST(\nRST~input_o ),
	.altera_internal_jtag1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

singlecycle CPU(
	.PC_29(\CPU|DP|PC [29]),
	.PC_28(\CPU|DP|PC [28]),
	.PC_31(\CPU|DP|PC [31]),
	.PC_30(\CPU|DP|PC [30]),
	.dpifhalt(\CPU|DP|dpif.halt~_Duplicate_1_q ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.LessThan1(\RAM|LessThan1~0_combout ),
	.PC_1(\CPU|DP|PC [1]),
	.daddr_1(\CPU|CM|daddr [1]),
	.ruifdWEN_r(\CPU|DP|ru|ruif.dWEN_r~q ),
	.ruifdREN_r(\CPU|DP|ru|ruif.dREN_r~q ),
	.daddr_0(\CPU|CM|daddr [0]),
	.PC_0(\CPU|DP|PC [0]),
	.daddr_3(\CPU|CM|daddr [3]),
	.PC_3(\CPU|DP|PC [3]),
	.daddr_2(\CPU|CM|daddr [2]),
	.PC_2(\CPU|DP|PC [2]),
	.daddr_5(\CPU|CM|daddr [5]),
	.PC_5(\CPU|DP|PC [5]),
	.daddr_4(\CPU|CM|daddr [4]),
	.PC_4(\CPU|DP|PC [4]),
	.daddr_7(\CPU|CM|daddr [7]),
	.PC_7(\CPU|DP|PC [7]),
	.daddr_6(\CPU|CM|daddr [6]),
	.PC_6(\CPU|DP|PC [6]),
	.always0(\RAM|always0~4_combout ),
	.daddr_9(\CPU|CM|daddr [9]),
	.PC_9(\CPU|DP|PC [9]),
	.PC_8(\CPU|DP|PC [8]),
	.daddr_8(\CPU|CM|daddr [8]),
	.daddr_11(\CPU|CM|daddr [11]),
	.PC_11(\CPU|DP|PC [11]),
	.daddr_10(\CPU|CM|daddr [10]),
	.PC_10(\CPU|DP|PC [10]),
	.daddr_13(\CPU|CM|daddr [13]),
	.PC_13(\CPU|DP|PC [13]),
	.daddr_12(\CPU|CM|daddr [12]),
	.PC_12(\CPU|DP|PC [12]),
	.daddr_15(\CPU|CM|daddr [15]),
	.PC_15(\CPU|DP|PC [15]),
	.daddr_14(\CPU|CM|daddr [14]),
	.PC_14(\CPU|DP|PC [14]),
	.always01(\RAM|always0~9_combout ),
	.PC_17(\CPU|DP|PC [17]),
	.daddr_17(\CPU|CM|daddr [17]),
	.daddr_16(\CPU|CM|daddr [16]),
	.PC_16(\CPU|DP|PC [16]),
	.daddr_19(\CPU|CM|daddr [19]),
	.PC_19(\CPU|DP|PC [19]),
	.daddr_18(\CPU|CM|daddr [18]),
	.PC_18(\CPU|DP|PC [18]),
	.PC_21(\CPU|DP|PC [21]),
	.daddr_21(\CPU|CM|daddr [21]),
	.PC_20(\CPU|DP|PC [20]),
	.daddr_20(\CPU|CM|daddr [20]),
	.daddr_23(\CPU|CM|daddr [23]),
	.PC_23(\CPU|DP|PC [23]),
	.daddr_22(\CPU|CM|daddr [22]),
	.PC_22(\CPU|DP|PC [22]),
	.daddr_25(\CPU|CM|daddr [25]),
	.PC_25(\CPU|DP|PC [25]),
	.daddr_24(\CPU|CM|daddr [24]),
	.PC_24(\CPU|DP|PC [24]),
	.daddr_27(\CPU|CM|daddr [27]),
	.PC_27(\CPU|DP|PC [27]),
	.daddr_26(\CPU|CM|daddr [26]),
	.PC_26(\CPU|DP|PC [26]),
	.daddr_29(\CPU|CM|daddr [29]),
	.daddr_28(\CPU|CM|daddr [28]),
	.daddr_31(\CPU|CM|daddr [31]),
	.daddr_30(\CPU|CM|daddr [30]),
	.always02(\RAM|always0~20_combout ),
	.always03(\RAM|always0~21_combout ),
	.ramiframload_01(\RAM|ramif.ramload[0]~1_combout ),
	.always1(\RAM|always1~1_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~2_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~3_combout ),
	.ramiframload_21(\RAM|ramif.ramload[2]~4_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~5_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~6_combout ),
	.ramiframload_41(\RAM|ramif.ramload[4]~7_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~8_combout ),
	.ramiframload_51(\RAM|ramif.ramload[5]~9_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~10_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~11_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~12_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~13_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~14_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~15_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~16_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~17_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~18_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~19_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~20_combout ),
	.ramiframload_161(\RAM|ramif.ramload[16]~21_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~22_combout ),
	.ramiframload_171(\RAM|ramif.ramload[17]~23_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~24_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~25_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~26_combout ),
	.ramiframload_211(\RAM|ramif.ramload[21]~27_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~28_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~29_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~30_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~31_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~32_combout ),
	.ramiframload_261(\RAM|ramif.ramload[26]~33_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~34_combout ),
	.ramiframload_271(\RAM|ramif.ramload[27]~35_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~36_combout ),
	.ramiframload_281(\RAM|ramif.ramload[28]~37_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~38_combout ),
	.ramiframload_291(\RAM|ramif.ramload[29]~39_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~40_combout ),
	.ramiframload_301(\RAM|ramif.ramload[30]~41_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~42_combout ),
	.ramiframload_311(\RAM|ramif.ramload[31]~43_combout ),
	.Mux63(\CPU|DP|rf|Mux63~9_combout ),
	.Mux631(\CPU|DP|rf|Mux63~19_combout ),
	.dcifimemload_20(\CPU|CM|dcif.imemload[20]~10_combout ),
	.Mux33(\CPU|DP|rf|Mux33~9_combout ),
	.Mux331(\CPU|DP|rf|Mux33~19_combout ),
	.Mux34(\CPU|DP|rf|Mux34~9_combout ),
	.Mux341(\CPU|DP|rf|Mux34~19_combout ),
	.Mux35(\CPU|DP|rf|Mux35~9_combout ),
	.Mux351(\CPU|DP|rf|Mux35~19_combout ),
	.Mux36(\CPU|DP|rf|Mux36~9_combout ),
	.Mux361(\CPU|DP|rf|Mux36~19_combout ),
	.Mux37(\CPU|DP|rf|Mux37~9_combout ),
	.Mux371(\CPU|DP|rf|Mux37~19_combout ),
	.Mux38(\CPU|DP|rf|Mux38~9_combout ),
	.Mux381(\CPU|DP|rf|Mux38~19_combout ),
	.Mux39(\CPU|DP|rf|Mux39~9_combout ),
	.Mux391(\CPU|DP|rf|Mux39~19_combout ),
	.Mux40(\CPU|DP|rf|Mux40~9_combout ),
	.Mux401(\CPU|DP|rf|Mux40~19_combout ),
	.Mux41(\CPU|DP|rf|Mux41~9_combout ),
	.Mux411(\CPU|DP|rf|Mux41~19_combout ),
	.Mux42(\CPU|DP|rf|Mux42~9_combout ),
	.Mux421(\CPU|DP|rf|Mux42~19_combout ),
	.Mux43(\CPU|DP|rf|Mux43~9_combout ),
	.Mux431(\CPU|DP|rf|Mux43~19_combout ),
	.Mux44(\CPU|DP|rf|Mux44~9_combout ),
	.Mux441(\CPU|DP|rf|Mux44~19_combout ),
	.Mux45(\CPU|DP|rf|Mux45~9_combout ),
	.Mux451(\CPU|DP|rf|Mux45~19_combout ),
	.Mux46(\CPU|DP|rf|Mux46~9_combout ),
	.Mux461(\CPU|DP|rf|Mux46~19_combout ),
	.Mux47(\CPU|DP|rf|Mux47~9_combout ),
	.Mux471(\CPU|DP|rf|Mux47~19_combout ),
	.Mux48(\CPU|DP|rf|Mux48~9_combout ),
	.Mux481(\CPU|DP|rf|Mux48~19_combout ),
	.Mux49(\CPU|DP|rf|Mux49~9_combout ),
	.Mux491(\CPU|DP|rf|Mux49~19_combout ),
	.Mux50(\CPU|DP|rf|Mux50~9_combout ),
	.Mux501(\CPU|DP|rf|Mux50~19_combout ),
	.Mux51(\CPU|DP|rf|Mux51~9_combout ),
	.Mux511(\CPU|DP|rf|Mux51~19_combout ),
	.Mux52(\CPU|DP|rf|Mux52~9_combout ),
	.Mux521(\CPU|DP|rf|Mux52~19_combout ),
	.Mux53(\CPU|DP|rf|Mux53~9_combout ),
	.Mux531(\CPU|DP|rf|Mux53~19_combout ),
	.Mux54(\CPU|DP|rf|Mux54~9_combout ),
	.Mux541(\CPU|DP|rf|Mux54~19_combout ),
	.Mux55(\CPU|DP|rf|Mux55~9_combout ),
	.Mux551(\CPU|DP|rf|Mux55~19_combout ),
	.Mux56(\CPU|DP|rf|Mux56~9_combout ),
	.Mux561(\CPU|DP|rf|Mux56~19_combout ),
	.Mux57(\CPU|DP|rf|Mux57~9_combout ),
	.Mux571(\CPU|DP|rf|Mux57~19_combout ),
	.Mux58(\CPU|DP|rf|Mux58~9_combout ),
	.Mux581(\CPU|DP|rf|Mux58~19_combout ),
	.Mux59(\CPU|DP|rf|Mux59~9_combout ),
	.Mux591(\CPU|DP|rf|Mux59~19_combout ),
	.Mux60(\CPU|DP|rf|Mux60~9_combout ),
	.Mux601(\CPU|DP|rf|Mux60~19_combout ),
	.Mux61(\CPU|DP|rf|Mux61~9_combout ),
	.Mux611(\CPU|DP|rf|Mux61~19_combout ),
	.Mux62(\CPU|DP|rf|Mux62~9_combout ),
	.Mux621(\CPU|DP|rf|Mux62~19_combout ),
	.Mux32(\CPU|DP|rf|Mux32~9_combout ),
	.Mux321(\CPU|DP|rf|Mux32~19_combout ),
	.nRST(\nRST~input_o ),
	.CLK(\CPUCLK~clkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.dpifhalt1(\CPU|DP|dpif.halt~q ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X56_Y37_N18
cycloneive_lcell_comb \ramaddr~0 (
// Equation(s):
// \ramaddr~0_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[1]~input_o )) # (!\syif.tbCTRL~input_o  & (((!ruifdREN_r & !ruifdWEN_r))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[1]~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~0 .lut_mask = 16'h888D;
defparam \ramaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N4
cycloneive_lcell_comb \ramaddr~1 (
// Equation(s):
// \ramaddr~1_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~0_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~0_combout  & (PC_1)) # (!\ramaddr~0_combout  & ((daddr_1)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC [1]),
	.datac(\CPU|CM|daddr [1]),
	.datad(\ramaddr~0_combout ),
	.cin(gnd),
	.combout(\ramaddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~1 .lut_mask = 16'hEE50;
defparam \ramaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N12
cycloneive_lcell_comb \ramaddr~2 (
// Equation(s):
// \ramaddr~2_combout  = (ruifdREN_r & (((daddr_0)))) # (!ruifdREN_r & ((ruifdWEN_r & ((daddr_0))) # (!ruifdWEN_r & (PC_0))))

	.dataa(\CPU|DP|ru|ruif.dREN_r~q ),
	.datab(\CPU|DP|PC [0]),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|CM|daddr [0]),
	.cin(gnd),
	.combout(\ramaddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~2 .lut_mask = 16'hFE04;
defparam \ramaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N6
cycloneive_lcell_comb \ramaddr~3 (
// Equation(s):
// \ramaddr~3_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~2_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[0]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~2_combout ),
	.cin(gnd),
	.combout(\ramaddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~3 .lut_mask = 16'hDD88;
defparam \ramaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N22
cycloneive_lcell_comb \ramaddr~4 (
// Equation(s):
// \ramaddr~4_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[3]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdREN_r) # (ruifdWEN_r))))

	.dataa(\syif.addr[3]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~4 .lut_mask = 16'hBBB8;
defparam \ramaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N26
cycloneive_lcell_comb \ramaddr~5 (
// Equation(s):
// \ramaddr~5_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~4_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~4_combout  & ((daddr_3))) # (!\ramaddr~4_combout  & (PC_3))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC [3]),
	.datac(\ramaddr~4_combout ),
	.datad(\CPU|CM|daddr [3]),
	.cin(gnd),
	.combout(\ramaddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~5 .lut_mask = 16'hF4A4;
defparam \ramaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N24
cycloneive_lcell_comb \ramaddr~6 (
// Equation(s):
// \ramaddr~6_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[2]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdREN_r) # (ruifdWEN_r))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[2]~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~6 .lut_mask = 16'hDDD8;
defparam \ramaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N2
cycloneive_lcell_comb \ramaddr~7 (
// Equation(s):
// \ramaddr~7_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~6_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~6_combout  & ((daddr_2))) # (!\ramaddr~6_combout  & (PC_2))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC [2]),
	.datac(\CPU|CM|daddr [2]),
	.datad(\ramaddr~6_combout ),
	.cin(gnd),
	.combout(\ramaddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~7 .lut_mask = 16'hFA44;
defparam \ramaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N16
cycloneive_lcell_comb \ramaddr~8 (
// Equation(s):
// \ramaddr~8_combout  = (ruifdREN_r & (((daddr_5)))) # (!ruifdREN_r & ((ruifdWEN_r & (daddr_5)) # (!ruifdWEN_r & ((PC_5)))))

	.dataa(\CPU|DP|ru|ruif.dREN_r~q ),
	.datab(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datac(\CPU|CM|daddr [5]),
	.datad(\CPU|DP|PC [5]),
	.cin(gnd),
	.combout(\ramaddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~8 .lut_mask = 16'hF1E0;
defparam \ramaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N2
cycloneive_lcell_comb \ramaddr~9 (
// Equation(s):
// \ramaddr~9_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~8_combout )))

	.dataa(\syif.addr[5]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~8_combout ),
	.cin(gnd),
	.combout(\ramaddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~9 .lut_mask = 16'hBB88;
defparam \ramaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N30
cycloneive_lcell_comb \ramaddr~10 (
// Equation(s):
// \ramaddr~10_combout  = (ruifdWEN_r & (((daddr_4)))) # (!ruifdWEN_r & ((ruifdREN_r & ((daddr_4))) # (!ruifdREN_r & (PC_4))))

	.dataa(\CPU|DP|PC [4]),
	.datab(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|CM|daddr [4]),
	.cin(gnd),
	.combout(\ramaddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~10 .lut_mask = 16'hFE02;
defparam \ramaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N20
cycloneive_lcell_comb \ramaddr~11 (
// Equation(s):
// \ramaddr~11_combout  = (\syif.tbCTRL~input_o  & ((\syif.addr[4]~input_o ))) # (!\syif.tbCTRL~input_o  & (\ramaddr~10_combout ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~10_combout ),
	.datad(\syif.addr[4]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~11 .lut_mask = 16'hFC30;
defparam \ramaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N2
cycloneive_lcell_comb \ramaddr~12 (
// Equation(s):
// \ramaddr~12_combout  = (ruifdWEN_r & (((daddr_7)))) # (!ruifdWEN_r & ((ruifdREN_r & ((daddr_7))) # (!ruifdREN_r & (PC_7))))

	.dataa(\CPU|DP|PC [7]),
	.datab(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|CM|daddr [7]),
	.cin(gnd),
	.combout(\ramaddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~12 .lut_mask = 16'hFE02;
defparam \ramaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N12
cycloneive_lcell_comb \ramaddr~13 (
// Equation(s):
// \ramaddr~13_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~12_combout )))

	.dataa(\syif.addr[7]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~12_combout ),
	.cin(gnd),
	.combout(\ramaddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~13 .lut_mask = 16'hAFA0;
defparam \ramaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N22
cycloneive_lcell_comb \ramaddr~14 (
// Equation(s):
// \ramaddr~14_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[6]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdWEN_r) # (ruifdREN_r))))

	.dataa(\syif.addr[6]~input_o ),
	.datab(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~14 .lut_mask = 16'hAAFC;
defparam \ramaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N24
cycloneive_lcell_comb \ramaddr~15 (
// Equation(s):
// \ramaddr~15_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~14_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~14_combout  & (daddr_6)) # (!\ramaddr~14_combout  & ((PC_6)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [6]),
	.datac(\ramaddr~14_combout ),
	.datad(\CPU|DP|PC [6]),
	.cin(gnd),
	.combout(\ramaddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~15 .lut_mask = 16'hE5E0;
defparam \ramaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N12
cycloneive_lcell_comb \ramaddr~16 (
// Equation(s):
// \ramaddr~16_combout  = (ruifdREN_r & (((daddr_9)))) # (!ruifdREN_r & ((ruifdWEN_r & ((daddr_9))) # (!ruifdWEN_r & (PC_9))))

	.dataa(\CPU|DP|PC [9]),
	.datab(\CPU|DP|ru|ruif.dREN_r~q ),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|CM|daddr [9]),
	.cin(gnd),
	.combout(\ramaddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~16 .lut_mask = 16'hFE02;
defparam \ramaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N18
cycloneive_lcell_comb \ramaddr~17 (
// Equation(s):
// \ramaddr~17_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~16_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[9]~input_o ),
	.datad(\ramaddr~16_combout ),
	.cin(gnd),
	.combout(\ramaddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~17 .lut_mask = 16'hF5A0;
defparam \ramaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N6
cycloneive_lcell_comb \ramaddr~18 (
// Equation(s):
// \ramaddr~18_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[8]~input_o )) # (!\syif.tbCTRL~input_o  & (((!ruifdWEN_r & !ruifdREN_r))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[8]~input_o ),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|DP|ru|ruif.dREN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~18 .lut_mask = 16'h888D;
defparam \ramaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N24
cycloneive_lcell_comb \ramaddr~19 (
// Equation(s):
// \ramaddr~19_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~18_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~18_combout  & (PC_8)) # (!\ramaddr~18_combout  & ((daddr_8)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC [8]),
	.datac(\CPU|CM|daddr [8]),
	.datad(\ramaddr~18_combout ),
	.cin(gnd),
	.combout(\ramaddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~19 .lut_mask = 16'hEE50;
defparam \ramaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N18
cycloneive_lcell_comb \ramaddr~20 (
// Equation(s):
// \ramaddr~20_combout  = (ruifdWEN_r & (((daddr_11)))) # (!ruifdWEN_r & ((ruifdREN_r & ((daddr_11))) # (!ruifdREN_r & (PC_11))))

	.dataa(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datab(\CPU|DP|PC [11]),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|CM|daddr [11]),
	.cin(gnd),
	.combout(\ramaddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~20 .lut_mask = 16'hFE04;
defparam \ramaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N12
cycloneive_lcell_comb \ramaddr~21 (
// Equation(s):
// \ramaddr~21_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~20_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[11]~input_o ),
	.datad(\ramaddr~20_combout ),
	.cin(gnd),
	.combout(\ramaddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~21 .lut_mask = 16'hF3C0;
defparam \ramaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N20
cycloneive_lcell_comb \ramaddr~22 (
// Equation(s):
// \ramaddr~22_combout  = (ruifdREN_r & (((daddr_10)))) # (!ruifdREN_r & ((ruifdWEN_r & ((daddr_10))) # (!ruifdWEN_r & (PC_10))))

	.dataa(\CPU|DP|PC [10]),
	.datab(\CPU|DP|ru|ruif.dREN_r~q ),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|CM|daddr [10]),
	.cin(gnd),
	.combout(\ramaddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~22 .lut_mask = 16'hFE02;
defparam \ramaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N10
cycloneive_lcell_comb \ramaddr~23 (
// Equation(s):
// \ramaddr~23_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~22_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[10]~input_o ),
	.datad(\ramaddr~22_combout ),
	.cin(gnd),
	.combout(\ramaddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~23 .lut_mask = 16'hF3C0;
defparam \ramaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N2
cycloneive_lcell_comb \ramaddr~24 (
// Equation(s):
// \ramaddr~24_combout  = (ruifdREN_r & (((daddr_13)))) # (!ruifdREN_r & ((ruifdWEN_r & ((daddr_13))) # (!ruifdWEN_r & (PC_13))))

	.dataa(\CPU|DP|PC [13]),
	.datab(\CPU|DP|ru|ruif.dREN_r~q ),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|CM|daddr [13]),
	.cin(gnd),
	.combout(\ramaddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~24 .lut_mask = 16'hFE02;
defparam \ramaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N16
cycloneive_lcell_comb \ramaddr~25 (
// Equation(s):
// \ramaddr~25_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[13]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~24_combout )))

	.dataa(gnd),
	.datab(\syif.addr[13]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~24_combout ),
	.cin(gnd),
	.combout(\ramaddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25 .lut_mask = 16'hCFC0;
defparam \ramaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N12
cycloneive_lcell_comb \ramaddr~26 (
// Equation(s):
// \ramaddr~26_combout  = (ruifdREN_r & (((daddr_12)))) # (!ruifdREN_r & ((ruifdWEN_r & ((daddr_12))) # (!ruifdWEN_r & (PC_12))))

	.dataa(\CPU|DP|PC [12]),
	.datab(\CPU|DP|ru|ruif.dREN_r~q ),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|CM|daddr [12]),
	.cin(gnd),
	.combout(\ramaddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~26 .lut_mask = 16'hFE02;
defparam \ramaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N18
cycloneive_lcell_comb \ramaddr~27 (
// Equation(s):
// \ramaddr~27_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~26_combout )))

	.dataa(gnd),
	.datab(\syif.addr[12]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~26_combout ),
	.cin(gnd),
	.combout(\ramaddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27 .lut_mask = 16'hCFC0;
defparam \ramaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N6
cycloneive_lcell_comb \ramaddr~28 (
// Equation(s):
// \ramaddr~28_combout  = (ruifdWEN_r & (((daddr_15)))) # (!ruifdWEN_r & ((ruifdREN_r & ((daddr_15))) # (!ruifdREN_r & (PC_15))))

	.dataa(\CPU|DP|PC [15]),
	.datab(\CPU|CM|daddr [15]),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|DP|ru|ruif.dREN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~28 .lut_mask = 16'hCCCA;
defparam \ramaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N24
cycloneive_lcell_comb \ramaddr~29 (
// Equation(s):
// \ramaddr~29_combout  = (\syif.tbCTRL~input_o  & (!\syif.addr[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~28_combout )))

	.dataa(\syif.addr[15]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~28_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29 .lut_mask = 16'h4477;
defparam \ramaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N0
cycloneive_lcell_comb \ramaddr~30 (
// Equation(s):
// \ramaddr~30_combout  = (ruifdWEN_r & (daddr_14)) # (!ruifdWEN_r & ((ruifdREN_r & (daddr_14)) # (!ruifdREN_r & ((PC_14)))))

	.dataa(\CPU|CM|daddr [14]),
	.datab(\CPU|DP|PC [14]),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|DP|ru|ruif.dREN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~30 .lut_mask = 16'hAAAC;
defparam \ramaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N2
cycloneive_lcell_comb \ramaddr~31 (
// Equation(s):
// \ramaddr~31_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~30_combout )))

	.dataa(\syif.addr[14]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~30_combout ),
	.cin(gnd),
	.combout(\ramaddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~31 .lut_mask = 16'hBB88;
defparam \ramaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N6
cycloneive_lcell_comb \ramaddr~32 (
// Equation(s):
// \ramaddr~32_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[17]~input_o )) # (!\syif.tbCTRL~input_o  & (((!ruifdREN_r & !ruifdWEN_r))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[17]~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~32 .lut_mask = 16'h888D;
defparam \ramaddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N16
cycloneive_lcell_comb \ramaddr~33 (
// Equation(s):
// \ramaddr~33_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~32_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~32_combout  & (PC_17)) # (!\ramaddr~32_combout  & ((daddr_17)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC [17]),
	.datac(\CPU|CM|daddr [17]),
	.datad(\ramaddr~32_combout ),
	.cin(gnd),
	.combout(\ramaddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~33 .lut_mask = 16'hEE50;
defparam \ramaddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N12
cycloneive_lcell_comb \ramaddr~34 (
// Equation(s):
// \ramaddr~34_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[16]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdREN_r) # (ruifdWEN_r))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[16]~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~34 .lut_mask = 16'hDDD8;
defparam \ramaddr~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N18
cycloneive_lcell_comb \ramaddr~35 (
// Equation(s):
// \ramaddr~35_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~34_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~34_combout  & (daddr_16)) # (!\ramaddr~34_combout  & ((PC_16)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [16]),
	.datac(\CPU|DP|PC [16]),
	.datad(\ramaddr~34_combout ),
	.cin(gnd),
	.combout(\ramaddr~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~35 .lut_mask = 16'hEE50;
defparam \ramaddr~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N10
cycloneive_lcell_comb \ramaddr~36 (
// Equation(s):
// \ramaddr~36_combout  = (ruifdREN_r & (daddr_19)) # (!ruifdREN_r & ((ruifdWEN_r & (daddr_19)) # (!ruifdWEN_r & ((PC_19)))))

	.dataa(\CPU|CM|daddr [19]),
	.datab(\CPU|DP|PC [19]),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~36 .lut_mask = 16'hAAAC;
defparam \ramaddr~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N6
cycloneive_lcell_comb \ramaddr~37 (
// Equation(s):
// \ramaddr~37_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~36_combout )))

	.dataa(\syif.addr[19]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~36_combout ),
	.cin(gnd),
	.combout(\ramaddr~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~37 .lut_mask = 16'hBB88;
defparam \ramaddr~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N18
cycloneive_lcell_comb \ramaddr~38 (
// Equation(s):
// \ramaddr~38_combout  = (ruifdWEN_r & (((daddr_18)))) # (!ruifdWEN_r & ((ruifdREN_r & ((daddr_18))) # (!ruifdREN_r & (PC_18))))

	.dataa(\CPU|DP|PC [18]),
	.datab(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|CM|daddr [18]),
	.cin(gnd),
	.combout(\ramaddr~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~38 .lut_mask = 16'hFE02;
defparam \ramaddr~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N16
cycloneive_lcell_comb \ramaddr~39 (
// Equation(s):
// \ramaddr~39_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~38_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[18]~input_o ),
	.datad(\ramaddr~38_combout ),
	.cin(gnd),
	.combout(\ramaddr~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~39 .lut_mask = 16'hF3C0;
defparam \ramaddr~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N30
cycloneive_lcell_comb \ramaddr~40 (
// Equation(s):
// \ramaddr~40_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[21]~input_o )))) # (!\syif.tbCTRL~input_o  & (!ruifdREN_r & ((!ruifdWEN_r))))

	.dataa(\CPU|DP|ru|ruif.dREN_r~q ),
	.datab(\syif.addr[21]~input_o ),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~40 .lut_mask = 16'hCC05;
defparam \ramaddr~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N24
cycloneive_lcell_comb \ramaddr~41 (
// Equation(s):
// \ramaddr~41_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~40_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~40_combout  & (PC_21)) # (!\ramaddr~40_combout  & ((daddr_21)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC [21]),
	.datac(\ramaddr~40_combout ),
	.datad(\CPU|CM|daddr [21]),
	.cin(gnd),
	.combout(\ramaddr~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~41 .lut_mask = 16'hE5E0;
defparam \ramaddr~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N20
cycloneive_lcell_comb \ramaddr~42 (
// Equation(s):
// \ramaddr~42_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[20]~input_o )))) # (!\syif.tbCTRL~input_o  & (!ruifdREN_r & ((!ruifdWEN_r))))

	.dataa(\CPU|DP|ru|ruif.dREN_r~q ),
	.datab(\syif.addr[20]~input_o ),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~42 .lut_mask = 16'hCC05;
defparam \ramaddr~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N18
cycloneive_lcell_comb \ramaddr~43 (
// Equation(s):
// \ramaddr~43_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~42_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~42_combout  & (PC_20)) # (!\ramaddr~42_combout  & ((daddr_20)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC [20]),
	.datac(\CPU|CM|daddr [20]),
	.datad(\ramaddr~42_combout ),
	.cin(gnd),
	.combout(\ramaddr~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~43 .lut_mask = 16'hEE50;
defparam \ramaddr~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N6
cycloneive_lcell_comb \ramaddr~44 (
// Equation(s):
// \ramaddr~44_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[23]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdREN_r) # (ruifdWEN_r))))

	.dataa(\syif.addr[23]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~44 .lut_mask = 16'hBBB8;
defparam \ramaddr~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N12
cycloneive_lcell_comb \ramaddr~45 (
// Equation(s):
// \ramaddr~45_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~44_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~44_combout  & (daddr_23)) # (!\ramaddr~44_combout  & ((PC_23)))))

	.dataa(\CPU|CM|daddr [23]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PC [23]),
	.datad(\ramaddr~44_combout ),
	.cin(gnd),
	.combout(\ramaddr~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~45 .lut_mask = 16'hEE30;
defparam \ramaddr~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N24
cycloneive_lcell_comb \ramaddr~46 (
// Equation(s):
// \ramaddr~46_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[22]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdREN_r) # (ruifdWEN_r))))

	.dataa(\syif.addr[22]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~46 .lut_mask = 16'hBBB8;
defparam \ramaddr~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N18
cycloneive_lcell_comb \ramaddr~47 (
// Equation(s):
// \ramaddr~47_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~46_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~46_combout  & ((daddr_22))) # (!\ramaddr~46_combout  & (PC_22))))

	.dataa(\CPU|DP|PC [22]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|daddr [22]),
	.datad(\ramaddr~46_combout ),
	.cin(gnd),
	.combout(\ramaddr~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~47 .lut_mask = 16'hFC22;
defparam \ramaddr~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N2
cycloneive_lcell_comb \ramaddr~48 (
// Equation(s):
// \ramaddr~48_combout  = (ruifdWEN_r & (((daddr_25)))) # (!ruifdWEN_r & ((ruifdREN_r & ((daddr_25))) # (!ruifdREN_r & (PC_25))))

	.dataa(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datab(\CPU|DP|PC [25]),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|CM|daddr [25]),
	.cin(gnd),
	.combout(\ramaddr~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~48 .lut_mask = 16'hFE04;
defparam \ramaddr~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N16
cycloneive_lcell_comb \ramaddr~49 (
// Equation(s):
// \ramaddr~49_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[25]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~48_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[25]~input_o ),
	.datad(\ramaddr~48_combout ),
	.cin(gnd),
	.combout(\ramaddr~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~49 .lut_mask = 16'hF3C0;
defparam \ramaddr~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N0
cycloneive_lcell_comb \ramaddr~50 (
// Equation(s):
// \ramaddr~50_combout  = (ruifdWEN_r & (((daddr_24)))) # (!ruifdWEN_r & ((ruifdREN_r & ((daddr_24))) # (!ruifdREN_r & (PC_24))))

	.dataa(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datab(\CPU|DP|ru|ruif.dREN_r~q ),
	.datac(\CPU|DP|PC [24]),
	.datad(\CPU|CM|daddr [24]),
	.cin(gnd),
	.combout(\ramaddr~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~50 .lut_mask = 16'hFE10;
defparam \ramaddr~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N30
cycloneive_lcell_comb \ramaddr~51 (
// Equation(s):
// \ramaddr~51_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~50_combout )))

	.dataa(gnd),
	.datab(\syif.addr[24]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~50_combout ),
	.cin(gnd),
	.combout(\ramaddr~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~51 .lut_mask = 16'hCFC0;
defparam \ramaddr~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N20
cycloneive_lcell_comb \ramaddr~52 (
// Equation(s):
// \ramaddr~52_combout  = (ruifdREN_r & (((daddr_27)))) # (!ruifdREN_r & ((ruifdWEN_r & ((daddr_27))) # (!ruifdWEN_r & (PC_27))))

	.dataa(\CPU|DP|ru|ruif.dREN_r~q ),
	.datab(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datac(\CPU|DP|PC [27]),
	.datad(\CPU|CM|daddr [27]),
	.cin(gnd),
	.combout(\ramaddr~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~52 .lut_mask = 16'hFE10;
defparam \ramaddr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N18
cycloneive_lcell_comb \ramaddr~53 (
// Equation(s):
// \ramaddr~53_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~52_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[27]~input_o ),
	.datad(\ramaddr~52_combout ),
	.cin(gnd),
	.combout(\ramaddr~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~53 .lut_mask = 16'hF5A0;
defparam \ramaddr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N2
cycloneive_lcell_comb \ramaddr~54 (
// Equation(s):
// \ramaddr~54_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[26]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdWEN_r) # (ruifdREN_r))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[26]~input_o ),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|DP|ru|ruif.dREN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~54 .lut_mask = 16'hDDD8;
defparam \ramaddr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N16
cycloneive_lcell_comb \ramaddr~55 (
// Equation(s):
// \ramaddr~55_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~54_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~54_combout  & (daddr_26)) # (!\ramaddr~54_combout  & ((PC_26)))))

	.dataa(\CPU|CM|daddr [26]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PC [26]),
	.datad(\ramaddr~54_combout ),
	.cin(gnd),
	.combout(\ramaddr~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~55 .lut_mask = 16'hEE30;
defparam \ramaddr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N6
cycloneive_lcell_comb \ramaddr~56 (
// Equation(s):
// \ramaddr~56_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[29]~input_o )) # (!\syif.tbCTRL~input_o  & (((!ruifdREN_r & !ruifdWEN_r))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[29]~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~56 .lut_mask = 16'h888D;
defparam \ramaddr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N20
cycloneive_lcell_comb \ramaddr~57 (
// Equation(s):
// \ramaddr~57_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~56_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~56_combout  & (PC_29)) # (!\ramaddr~56_combout  & ((daddr_29)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC [29]),
	.datac(\CPU|CM|daddr [29]),
	.datad(\ramaddr~56_combout ),
	.cin(gnd),
	.combout(\ramaddr~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~57 .lut_mask = 16'hEE50;
defparam \ramaddr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N28
cycloneive_lcell_comb \ramaddr~58 (
// Equation(s):
// \ramaddr~58_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[28]~input_o )) # (!\syif.tbCTRL~input_o  & (((!ruifdREN_r & !ruifdWEN_r))))

	.dataa(\syif.addr[28]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\CPU|DP|ru|ruif.dWEN_r~q ),
	.cin(gnd),
	.combout(\ramaddr~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~58 .lut_mask = 16'h888B;
defparam \ramaddr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N18
cycloneive_lcell_comb \ramaddr~59 (
// Equation(s):
// \ramaddr~59_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~58_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~58_combout  & (PC_28)) # (!\ramaddr~58_combout  & ((daddr_28)))))

	.dataa(\CPU|DP|PC [28]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|daddr [28]),
	.datad(\ramaddr~58_combout ),
	.cin(gnd),
	.combout(\ramaddr~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~59 .lut_mask = 16'hEE30;
defparam \ramaddr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N10
cycloneive_lcell_comb \ramaddr~60 (
// Equation(s):
// \ramaddr~60_combout  = (ruifdREN_r & (((daddr_31)))) # (!ruifdREN_r & ((ruifdWEN_r & ((daddr_31))) # (!ruifdWEN_r & (PC_31))))

	.dataa(\CPU|DP|ru|ruif.dREN_r~q ),
	.datab(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datac(\CPU|DP|PC [31]),
	.datad(\CPU|CM|daddr [31]),
	.cin(gnd),
	.combout(\ramaddr~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~60 .lut_mask = 16'hFE10;
defparam \ramaddr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N12
cycloneive_lcell_comb \ramaddr~61 (
// Equation(s):
// \ramaddr~61_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~60_combout )))

	.dataa(\syif.addr[31]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~60_combout ),
	.cin(gnd),
	.combout(\ramaddr~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~61 .lut_mask = 16'hAFA0;
defparam \ramaddr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N4
cycloneive_lcell_comb \ramaddr~62 (
// Equation(s):
// \ramaddr~62_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[30]~input_o )))) # (!\syif.tbCTRL~input_o  & ((ruifdREN_r) # ((ruifdWEN_r))))

	.dataa(\CPU|DP|ru|ruif.dREN_r~q ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\syif.addr[30]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~62 .lut_mask = 16'hFE32;
defparam \ramaddr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N18
cycloneive_lcell_comb \ramaddr~63 (
// Equation(s):
// \ramaddr~63_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~62_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~62_combout  & ((daddr_30))) # (!\ramaddr~62_combout  & (PC_30))))

	.dataa(\CPU|DP|PC [30]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~62_combout ),
	.datad(\CPU|CM|daddr [30]),
	.cin(gnd),
	.combout(\ramaddr~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~63 .lut_mask = 16'hF2C2;
defparam \ramaddr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N28
cycloneive_lcell_comb \ramWEN~0 (
// Equation(s):
// \ramWEN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.WEN~input_o )) # (!\syif.tbCTRL~input_o  & ((!ruifdWEN_r)))

	.dataa(\syif.WEN~input_o ),
	.datab(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~0 .lut_mask = 16'h5353;
defparam \ramWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N14
cycloneive_lcell_comb \ramREN~0 (
// Equation(s):
// \ramREN~0_combout  = (!\syif.tbCTRL~input_o  & (!ruifdWEN_r & !dpifhalt))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\CPU|DP|ru|ruif.dWEN_r~q ),
	.datad(\CPU|DP|dpif.halt~_Duplicate_1_q ),
	.cin(gnd),
	.combout(\ramREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~0 .lut_mask = 16'h0005;
defparam \ramREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N6
cycloneive_lcell_comb \ramREN~1 (
// Equation(s):
// \ramREN~1_combout  = (!\ramREN~0_combout  & ((\syif.tbCTRL~input_o  & (!\syif.REN~input_o )) # (!\syif.tbCTRL~input_o  & ((!ruifdREN_r)))))

	.dataa(\syif.REN~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru|ruif.dREN_r~q ),
	.datad(\ramREN~0_combout ),
	.cin(gnd),
	.combout(\ramREN~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~1 .lut_mask = 16'h0047;
defparam \ramREN~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X114_Y37_N17
dffeas CPUCLK(
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\CPUCLK~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\CPUCLK~q ),
	.prn(vcc));
// synopsys translate_off
defparam CPUCLK.is_wysiwyg = "true";
defparam CPUCLK.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N18
cycloneive_lcell_comb \ramstore~0 (
// Equation(s):
// \ramstore~0_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux63)) # (!dcifimemload_20 & ((Mux631)))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\CPU|DP|rf|Mux63~9_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf|Mux63~19_combout ),
	.cin(gnd),
	.combout(\ramstore~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~0 .lut_mask = 16'h0D08;
defparam \ramstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N4
cycloneive_lcell_comb \ramstore~1 (
// Equation(s):
// \ramstore~1_combout  = (\ramstore~0_combout ) # ((\syif.store[0]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[0]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~0_combout ),
	.cin(gnd),
	.combout(\ramstore~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~1 .lut_mask = 16'hFFC0;
defparam \ramstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N10
cycloneive_lcell_comb \ramstore~2 (
// Equation(s):
// \ramstore~2_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux62)) # (!dcifimemload_20 & ((Mux621)))))

	.dataa(\CPU|DP|rf|Mux62~9_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|rf|Mux62~19_combout ),
	.cin(gnd),
	.combout(\ramstore~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~2 .lut_mask = 16'h2320;
defparam \ramstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N16
cycloneive_lcell_comb \ramstore~3 (
// Equation(s):
// \ramstore~3_combout  = (\ramstore~2_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[1]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[1]~input_o ),
	.datad(\ramstore~2_combout ),
	.cin(gnd),
	.combout(\ramstore~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~3 .lut_mask = 16'hFFC0;
defparam \ramstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N2
cycloneive_lcell_comb \ramstore~4 (
// Equation(s):
// \ramstore~4_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux61)) # (!dcifimemload_20 & ((Mux611)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|rf|Mux61~9_combout ),
	.datad(\CPU|DP|rf|Mux61~19_combout ),
	.cin(gnd),
	.combout(\ramstore~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~4 .lut_mask = 16'h5140;
defparam \ramstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N4
cycloneive_lcell_comb \ramstore~5 (
// Equation(s):
// \ramstore~5_combout  = (\ramstore~4_combout ) # ((\syif.store[2]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[2]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~4_combout ),
	.cin(gnd),
	.combout(\ramstore~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~5 .lut_mask = 16'hFFC0;
defparam \ramstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N16
cycloneive_lcell_comb \ramstore~6 (
// Equation(s):
// \ramstore~6_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux60)) # (!dcifimemload_20 & ((Mux601)))))

	.dataa(\CPU|DP|rf|Mux60~9_combout ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf|Mux60~19_combout ),
	.cin(gnd),
	.combout(\ramstore~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~6 .lut_mask = 16'h0B08;
defparam \ramstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N14
cycloneive_lcell_comb \ramstore~7 (
// Equation(s):
// \ramstore~7_combout  = (\ramstore~6_combout ) # ((\syif.store[3]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[3]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~6_combout ),
	.cin(gnd),
	.combout(\ramstore~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~7 .lut_mask = 16'hFFA0;
defparam \ramstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N8
cycloneive_lcell_comb \ramstore~8 (
// Equation(s):
// \ramstore~8_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux59)) # (!dcifimemload_20 & ((Mux591)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|rf|Mux59~9_combout ),
	.datad(\CPU|DP|rf|Mux59~19_combout ),
	.cin(gnd),
	.combout(\ramstore~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~8 .lut_mask = 16'h5140;
defparam \ramstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N10
cycloneive_lcell_comb \ramstore~9 (
// Equation(s):
// \ramstore~9_combout  = (\ramstore~8_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[4]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[4]~input_o ),
	.datac(\ramstore~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~9 .lut_mask = 16'hF8F8;
defparam \ramstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N6
cycloneive_lcell_comb \ramstore~10 (
// Equation(s):
// \ramstore~10_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux58)) # (!dcifimemload_20 & ((Mux581)))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux58~9_combout ),
	.datad(\CPU|DP|rf|Mux58~19_combout ),
	.cin(gnd),
	.combout(\ramstore~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~10 .lut_mask = 16'h3120;
defparam \ramstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N0
cycloneive_lcell_comb \ramstore~11 (
// Equation(s):
// \ramstore~11_combout  = (\ramstore~10_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[5]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[5]~input_o ),
	.datad(\ramstore~10_combout ),
	.cin(gnd),
	.combout(\ramstore~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~11 .lut_mask = 16'hFFC0;
defparam \ramstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N0
cycloneive_lcell_comb \ramstore~12 (
// Equation(s):
// \ramstore~12_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux57))) # (!dcifimemload_20 & (Mux571))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux57~19_combout ),
	.datad(\CPU|DP|rf|Mux57~9_combout ),
	.cin(gnd),
	.combout(\ramstore~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~12 .lut_mask = 16'h3210;
defparam \ramstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N30
cycloneive_lcell_comb \ramstore~13 (
// Equation(s):
// \ramstore~13_combout  = (\ramstore~12_combout ) # ((\syif.store[6]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[6]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~12_combout ),
	.cin(gnd),
	.combout(\ramstore~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~13 .lut_mask = 16'hFFC0;
defparam \ramstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N20
cycloneive_lcell_comb \ramstore~14 (
// Equation(s):
// \ramstore~14_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux56)) # (!dcifimemload_20 & ((Mux561)))))

	.dataa(\CPU|DP|rf|Mux56~9_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|rf|Mux56~19_combout ),
	.cin(gnd),
	.combout(\ramstore~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~14 .lut_mask = 16'h2320;
defparam \ramstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N26
cycloneive_lcell_comb \ramstore~15 (
// Equation(s):
// \ramstore~15_combout  = (\ramstore~14_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[7]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[7]~input_o ),
	.datad(\ramstore~14_combout ),
	.cin(gnd),
	.combout(\ramstore~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~15 .lut_mask = 16'hFFC0;
defparam \ramstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N20
cycloneive_lcell_comb \ramstore~16 (
// Equation(s):
// \ramstore~16_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux55)) # (!dcifimemload_20 & ((Mux551)))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux55~9_combout ),
	.datad(\CPU|DP|rf|Mux55~19_combout ),
	.cin(gnd),
	.combout(\ramstore~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~16 .lut_mask = 16'h3120;
defparam \ramstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N18
cycloneive_lcell_comb \ramstore~17 (
// Equation(s):
// \ramstore~17_combout  = (\ramstore~16_combout ) # ((\syif.store[8]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[8]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~16_combout ),
	.cin(gnd),
	.combout(\ramstore~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~17 .lut_mask = 16'hFFA0;
defparam \ramstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N0
cycloneive_lcell_comb \ramstore~18 (
// Equation(s):
// \ramstore~18_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux54))) # (!dcifimemload_20 & (Mux541))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|rf|Mux54~19_combout ),
	.datad(\CPU|DP|rf|Mux54~9_combout ),
	.cin(gnd),
	.combout(\ramstore~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~18 .lut_mask = 16'h5410;
defparam \ramstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N22
cycloneive_lcell_comb \ramstore~19 (
// Equation(s):
// \ramstore~19_combout  = (\ramstore~18_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[9]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[9]~input_o ),
	.datad(\ramstore~18_combout ),
	.cin(gnd),
	.combout(\ramstore~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~19 .lut_mask = 16'hFFC0;
defparam \ramstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N12
cycloneive_lcell_comb \ramstore~20 (
// Equation(s):
// \ramstore~20_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux53))) # (!dcifimemload_20 & (Mux531))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux53~19_combout ),
	.datad(\CPU|DP|rf|Mux53~9_combout ),
	.cin(gnd),
	.combout(\ramstore~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~20 .lut_mask = 16'h3210;
defparam \ramstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N26
cycloneive_lcell_comb \ramstore~21 (
// Equation(s):
// \ramstore~21_combout  = (\ramstore~20_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[10]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[10]~input_o ),
	.datad(\ramstore~20_combout ),
	.cin(gnd),
	.combout(\ramstore~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~21 .lut_mask = 16'hFFC0;
defparam \ramstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N20
cycloneive_lcell_comb \ramstore~22 (
// Equation(s):
// \ramstore~22_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux52))) # (!dcifimemload_20 & (Mux521))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux52~19_combout ),
	.datad(\CPU|DP|rf|Mux52~9_combout ),
	.cin(gnd),
	.combout(\ramstore~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~22 .lut_mask = 16'h3210;
defparam \ramstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N10
cycloneive_lcell_comb \ramstore~23 (
// Equation(s):
// \ramstore~23_combout  = (\ramstore~22_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[11]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[11]~input_o ),
	.datad(\ramstore~22_combout ),
	.cin(gnd),
	.combout(\ramstore~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~23 .lut_mask = 16'hFFC0;
defparam \ramstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N20
cycloneive_lcell_comb \ramstore~24 (
// Equation(s):
// \ramstore~24_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux51)) # (!dcifimemload_20 & ((Mux511)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|rf|Mux51~9_combout ),
	.datad(\CPU|DP|rf|Mux51~19_combout ),
	.cin(gnd),
	.combout(\ramstore~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~24 .lut_mask = 16'h5140;
defparam \ramstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N14
cycloneive_lcell_comb \ramstore~25 (
// Equation(s):
// \ramstore~25_combout  = (\ramstore~24_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[12]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[12]~input_o ),
	.datac(gnd),
	.datad(\ramstore~24_combout ),
	.cin(gnd),
	.combout(\ramstore~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~25 .lut_mask = 16'hFF88;
defparam \ramstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N24
cycloneive_lcell_comb \ramstore~26 (
// Equation(s):
// \ramstore~26_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux50))) # (!dcifimemload_20 & (Mux501))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux50~19_combout ),
	.datad(\CPU|DP|rf|Mux50~9_combout ),
	.cin(gnd),
	.combout(\ramstore~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~26 .lut_mask = 16'h3210;
defparam \ramstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N6
cycloneive_lcell_comb \ramstore~27 (
// Equation(s):
// \ramstore~27_combout  = (\ramstore~26_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[13]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[13]~input_o ),
	.datad(\ramstore~26_combout ),
	.cin(gnd),
	.combout(\ramstore~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~27 .lut_mask = 16'hFFC0;
defparam \ramstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N28
cycloneive_lcell_comb \ramstore~28 (
// Equation(s):
// \ramstore~28_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux49))) # (!dcifimemload_20 & (Mux491))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux49~19_combout ),
	.datad(\CPU|DP|rf|Mux49~9_combout ),
	.cin(gnd),
	.combout(\ramstore~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~28 .lut_mask = 16'h3210;
defparam \ramstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N2
cycloneive_lcell_comb \ramstore~29 (
// Equation(s):
// \ramstore~29_combout  = (\ramstore~28_combout ) # ((\syif.store[14]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[14]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~28_combout ),
	.cin(gnd),
	.combout(\ramstore~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~29 .lut_mask = 16'hFFA0;
defparam \ramstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N6
cycloneive_lcell_comb \ramstore~30 (
// Equation(s):
// \ramstore~30_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux48))) # (!dcifimemload_20 & (Mux481))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux48~19_combout ),
	.datad(\CPU|DP|rf|Mux48~9_combout ),
	.cin(gnd),
	.combout(\ramstore~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~30 .lut_mask = 16'h3210;
defparam \ramstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N20
cycloneive_lcell_comb \ramstore~31 (
// Equation(s):
// \ramstore~31_combout  = (\ramstore~30_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[15]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[15]~input_o ),
	.datad(\ramstore~30_combout ),
	.cin(gnd),
	.combout(\ramstore~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~31 .lut_mask = 16'hFFC0;
defparam \ramstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N2
cycloneive_lcell_comb \ramstore~32 (
// Equation(s):
// \ramstore~32_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux47))) # (!dcifimemload_20 & (Mux471))))

	.dataa(\CPU|DP|rf|Mux47~19_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|rf|Mux47~9_combout ),
	.cin(gnd),
	.combout(\ramstore~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~32 .lut_mask = 16'h3202;
defparam \ramstore~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N28
cycloneive_lcell_comb \ramstore~33 (
// Equation(s):
// \ramstore~33_combout  = (\ramstore~32_combout ) # ((\syif.store[16]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[16]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramstore~32_combout ),
	.cin(gnd),
	.combout(\ramstore~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~33 .lut_mask = 16'hFF88;
defparam \ramstore~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N20
cycloneive_lcell_comb \ramstore~34 (
// Equation(s):
// \ramstore~34_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux46))) # (!dcifimemload_20 & (Mux461))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|rf|Mux46~19_combout ),
	.datad(\CPU|DP|rf|Mux46~9_combout ),
	.cin(gnd),
	.combout(\ramstore~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~34 .lut_mask = 16'h5410;
defparam \ramstore~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N14
cycloneive_lcell_comb \ramstore~35 (
// Equation(s):
// \ramstore~35_combout  = (\ramstore~34_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[17]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[17]~input_o ),
	.datad(\ramstore~34_combout ),
	.cin(gnd),
	.combout(\ramstore~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~35 .lut_mask = 16'hFFA0;
defparam \ramstore~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N20
cycloneive_lcell_comb \ramstore~36 (
// Equation(s):
// \ramstore~36_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux45))) # (!dcifimemload_20 & (Mux451))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\CPU|DP|rf|Mux45~19_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf|Mux45~9_combout ),
	.cin(gnd),
	.combout(\ramstore~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~36 .lut_mask = 16'h0E04;
defparam \ramstore~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N22
cycloneive_lcell_comb \ramstore~37 (
// Equation(s):
// \ramstore~37_combout  = (\ramstore~36_combout ) # ((\syif.store[18]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[18]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~36_combout ),
	.cin(gnd),
	.combout(\ramstore~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~37 .lut_mask = 16'hFFC0;
defparam \ramstore~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N20
cycloneive_lcell_comb \ramstore~38 (
// Equation(s):
// \ramstore~38_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux44))) # (!dcifimemload_20 & (Mux441))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\CPU|DP|rf|Mux44~19_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf|Mux44~9_combout ),
	.cin(gnd),
	.combout(\ramstore~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~38 .lut_mask = 16'h0E04;
defparam \ramstore~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N10
cycloneive_lcell_comb \ramstore~39 (
// Equation(s):
// \ramstore~39_combout  = (\ramstore~38_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[19]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[19]~input_o ),
	.datad(\ramstore~38_combout ),
	.cin(gnd),
	.combout(\ramstore~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~39 .lut_mask = 16'hFFC0;
defparam \ramstore~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N12
cycloneive_lcell_comb \ramstore~40 (
// Equation(s):
// \ramstore~40_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux43)) # (!dcifimemload_20 & ((Mux431)))))

	.dataa(\CPU|DP|rf|Mux43~9_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|rf|Mux43~19_combout ),
	.cin(gnd),
	.combout(\ramstore~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~40 .lut_mask = 16'h2320;
defparam \ramstore~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N18
cycloneive_lcell_comb \ramstore~41 (
// Equation(s):
// \ramstore~41_combout  = (\ramstore~40_combout ) # ((\syif.store[20]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[20]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~40_combout ),
	.cin(gnd),
	.combout(\ramstore~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~41 .lut_mask = 16'hFFC0;
defparam \ramstore~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N18
cycloneive_lcell_comb \ramstore~42 (
// Equation(s):
// \ramstore~42_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux42))) # (!dcifimemload_20 & (Mux421))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\CPU|DP|rf|Mux42~19_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf|Mux42~9_combout ),
	.cin(gnd),
	.combout(\ramstore~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~42 .lut_mask = 16'h0E04;
defparam \ramstore~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N0
cycloneive_lcell_comb \ramstore~43 (
// Equation(s):
// \ramstore~43_combout  = (\ramstore~42_combout ) # ((\syif.store[21]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[21]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~42_combout ),
	.cin(gnd),
	.combout(\ramstore~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~43 .lut_mask = 16'hFFC0;
defparam \ramstore~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N12
cycloneive_lcell_comb \ramstore~44 (
// Equation(s):
// \ramstore~44_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux41))) # (!dcifimemload_20 & (Mux411))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\CPU|DP|rf|Mux41~19_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf|Mux41~9_combout ),
	.cin(gnd),
	.combout(\ramstore~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~44 .lut_mask = 16'h0E04;
defparam \ramstore~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N22
cycloneive_lcell_comb \ramstore~45 (
// Equation(s):
// \ramstore~45_combout  = (\ramstore~44_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[22]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[22]~input_o ),
	.datad(\ramstore~44_combout ),
	.cin(gnd),
	.combout(\ramstore~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~45 .lut_mask = 16'hFFC0;
defparam \ramstore~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N24
cycloneive_lcell_comb \ramstore~46 (
// Equation(s):
// \ramstore~46_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux40))) # (!dcifimemload_20 & (Mux401))))

	.dataa(\CPU|DP|rf|Mux40~19_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux40~9_combout ),
	.datad(\CPU|CM|dcif.imemload[20]~10_combout ),
	.cin(gnd),
	.combout(\ramstore~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~46 .lut_mask = 16'h3022;
defparam \ramstore~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N14
cycloneive_lcell_comb \ramstore~47 (
// Equation(s):
// \ramstore~47_combout  = (\ramstore~46_combout ) # ((\syif.store[23]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[23]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramstore~46_combout ),
	.cin(gnd),
	.combout(\ramstore~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~47 .lut_mask = 16'hFF88;
defparam \ramstore~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N12
cycloneive_lcell_comb \ramstore~48 (
// Equation(s):
// \ramstore~48_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux39))) # (!dcifimemload_20 & (Mux391))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|rf|Mux39~19_combout ),
	.datad(\CPU|DP|rf|Mux39~9_combout ),
	.cin(gnd),
	.combout(\ramstore~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~48 .lut_mask = 16'h5410;
defparam \ramstore~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N22
cycloneive_lcell_comb \ramstore~49 (
// Equation(s):
// \ramstore~49_combout  = (\ramstore~48_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[24]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[24]~input_o ),
	.datad(\ramstore~48_combout ),
	.cin(gnd),
	.combout(\ramstore~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~49 .lut_mask = 16'hFFC0;
defparam \ramstore~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N28
cycloneive_lcell_comb \ramstore~50 (
// Equation(s):
// \ramstore~50_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux38))) # (!dcifimemload_20 & (Mux381))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux38~19_combout ),
	.datad(\CPU|DP|rf|Mux38~9_combout ),
	.cin(gnd),
	.combout(\ramstore~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~50 .lut_mask = 16'h3210;
defparam \ramstore~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N10
cycloneive_lcell_comb \ramstore~51 (
// Equation(s):
// \ramstore~51_combout  = (\ramstore~50_combout ) # ((\syif.store[25]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[25]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~50_combout ),
	.cin(gnd),
	.combout(\ramstore~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~51 .lut_mask = 16'hFFA0;
defparam \ramstore~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N24
cycloneive_lcell_comb \ramstore~52 (
// Equation(s):
// \ramstore~52_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux37))) # (!dcifimemload_20 & (Mux371))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|rf|Mux37~19_combout ),
	.datad(\CPU|DP|rf|Mux37~9_combout ),
	.cin(gnd),
	.combout(\ramstore~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~52 .lut_mask = 16'h5410;
defparam \ramstore~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N6
cycloneive_lcell_comb \ramstore~53 (
// Equation(s):
// \ramstore~53_combout  = (\ramstore~52_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[26]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[26]~input_o ),
	.datad(\ramstore~52_combout ),
	.cin(gnd),
	.combout(\ramstore~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~53 .lut_mask = 16'hFFA0;
defparam \ramstore~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N16
cycloneive_lcell_comb \ramstore~54 (
// Equation(s):
// \ramstore~54_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux36))) # (!dcifimemload_20 & (Mux361))))

	.dataa(\CPU|DP|rf|Mux36~19_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|rf|Mux36~9_combout ),
	.cin(gnd),
	.combout(\ramstore~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~54 .lut_mask = 16'h3202;
defparam \ramstore~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N22
cycloneive_lcell_comb \ramstore~55 (
// Equation(s):
// \ramstore~55_combout  = (\ramstore~54_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[27]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[27]~input_o ),
	.datad(\ramstore~54_combout ),
	.cin(gnd),
	.combout(\ramstore~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~55 .lut_mask = 16'hFFC0;
defparam \ramstore~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N12
cycloneive_lcell_comb \ramstore~56 (
// Equation(s):
// \ramstore~56_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux35)) # (!dcifimemload_20 & ((Mux351)))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux35~9_combout ),
	.datad(\CPU|DP|rf|Mux35~19_combout ),
	.cin(gnd),
	.combout(\ramstore~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~56 .lut_mask = 16'h3120;
defparam \ramstore~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N14
cycloneive_lcell_comb \ramstore~57 (
// Equation(s):
// \ramstore~57_combout  = (\ramstore~56_combout ) # ((\syif.store[28]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[28]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~56_combout ),
	.cin(gnd),
	.combout(\ramstore~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~57 .lut_mask = 16'hFFA0;
defparam \ramstore~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N28
cycloneive_lcell_comb \ramstore~58 (
// Equation(s):
// \ramstore~58_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux34))) # (!dcifimemload_20 & (Mux341))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|rf|Mux34~19_combout ),
	.datad(\CPU|DP|rf|Mux34~9_combout ),
	.cin(gnd),
	.combout(\ramstore~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~58 .lut_mask = 16'h5410;
defparam \ramstore~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N26
cycloneive_lcell_comb \ramstore~59 (
// Equation(s):
// \ramstore~59_combout  = (\ramstore~58_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[29]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[29]~input_o ),
	.datad(\ramstore~58_combout ),
	.cin(gnd),
	.combout(\ramstore~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~59 .lut_mask = 16'hFFC0;
defparam \ramstore~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N28
cycloneive_lcell_comb \ramstore~60 (
// Equation(s):
// \ramstore~60_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux33))) # (!dcifimemload_20 & (Mux331))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf|Mux33~19_combout ),
	.datad(\CPU|DP|rf|Mux33~9_combout ),
	.cin(gnd),
	.combout(\ramstore~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~60 .lut_mask = 16'h3210;
defparam \ramstore~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N2
cycloneive_lcell_comb \ramstore~61 (
// Equation(s):
// \ramstore~61_combout  = (\ramstore~60_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[30]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[30]~input_o ),
	.datad(\ramstore~60_combout ),
	.cin(gnd),
	.combout(\ramstore~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~61 .lut_mask = 16'hFFC0;
defparam \ramstore~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N28
cycloneive_lcell_comb \ramstore~62 (
// Equation(s):
// \ramstore~62_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux321))) # (!dcifimemload_20 & (Mux32))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\CPU|DP|rf|Mux32~9_combout ),
	.datac(\CPU|DP|rf|Mux32~19_combout ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~62 .lut_mask = 16'h00E4;
defparam \ramstore~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N22
cycloneive_lcell_comb \ramstore~63 (
// Equation(s):
// \ramstore~63_combout  = (\ramstore~62_combout ) # ((\syif.store[31]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[31]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~62_combout ),
	.cin(gnd),
	.combout(\ramstore~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~63 .lut_mask = 16'hFFC0;
defparam \ramstore~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X113_Y37_N1
dffeas \count[3] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X113_Y37_N23
dffeas \count[2] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X113_Y37_N13
dffeas \count[1] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X113_Y37_N3
dffeas \count[0] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X113_Y37_N24
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!count[1] & (!count[0] & (!count[2] & !count[3])))

	.dataa(count[1]),
	.datab(count[0]),
	.datac(count[2]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X114_Y37_N16
cycloneive_lcell_comb \CPUCLK~0 (
// Equation(s):
// \CPUCLK~0_combout  = \CPUCLK~q  $ (\Equal0~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\CPUCLK~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\CPUCLK~0_combout ),
	.cout());
// synopsys translate_off
defparam \CPUCLK~0 .lut_mask = 16'h0FF0;
defparam \CPUCLK~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X113_Y37_N0
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = count[3] $ (((count[2] & (count[0] & count[1]))))

	.dataa(count[2]),
	.datab(count[0]),
	.datac(count[3]),
	.datad(count[1]),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h78F0;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X113_Y37_N22
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = count[2] $ (((count[0] & count[1])))

	.dataa(gnd),
	.datab(count[0]),
	.datac(count[2]),
	.datad(count[1]),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h3CF0;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X113_Y37_N12
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = count[1] $ (count[0])

	.dataa(gnd),
	.datab(gnd),
	.datac(count[1]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h0FF0;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X113_Y37_N2
cycloneive_lcell_comb \count~3 (
// Equation(s):
// \count~3_combout  = (!count[0] & ((count[2]) # ((count[3]) # (count[1]))))

	.dataa(count[2]),
	.datab(count[3]),
	.datac(count[0]),
	.datad(count[1]),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
// synopsys translate_off
defparam \count~3 .lut_mask = 16'h0F0E;
defparam \count~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N26
cycloneive_lcell_comb \ramaddr~29_wirecell (
// Equation(s):
// \ramaddr~29_wirecell_combout  = !\ramaddr~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\ramaddr~29_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29_wirecell .lut_mask = 16'h00FF;
defparam \ramaddr~29_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: JTAG_X1_Y37_N0
cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

// Location: FF_X43_Y39_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y36_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y39_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .lut_mask = 16'hEE44;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y36_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y39_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~10 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~10 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 .lut_mask = 16'h5AAF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .lut_mask = 16'h5A5A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y36_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hC30C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .lut_mask = 16'hA5A5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .lut_mask = 16'h33AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y36_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .lut_mask = 16'hDD88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y39_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .lut_mask = 16'hF870;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .lut_mask = 16'h004C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .lut_mask = 16'hF0A8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .lut_mask = 16'h88B8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 .lut_mask = 16'h0003;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5 .lut_mask = 16'h43C4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .lut_mask = 16'hC0F3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7 .lut_mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .lut_mask = 16'h00F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .lut_mask = 16'h33FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .lut_mask = 16'hFC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .lut_mask = 16'h8081;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y38_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .lut_mask = 16'hCECC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .lut_mask = 16'h0C0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .lut_mask = 16'h5C02;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .lut_mask = 16'hD2F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .lut_mask = 16'h0080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y39_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .lut_mask = 16'h5AF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7 .lut_mask = 16'hFF04;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8 .lut_mask = 16'hF888;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .lut_mask = 16'h0200;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .lut_mask = 16'hDADA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .lut_mask = 16'hCECE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .lut_mask = 16'h4121;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y38_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .lut_mask = 16'h8D88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .lut_mask = 16'h0C0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y36_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .lut_mask = 16'h2200;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .lut_mask = 16'h8B26;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .lut_mask = 16'hC0F3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .lut_mask = 16'hAAAB;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .lut_mask = 16'h0100;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y38_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .lut_mask = 16'hCECC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y36_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .lut_mask = 16'h0030;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .lut_mask = 16'hD407;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .lut_mask = 16'hF3C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .lut_mask = 16'h1110;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .lut_mask = 16'h0E0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y36_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .lut_mask = 16'hFFC8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hCE0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hFF40;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .lut_mask = 16'h2A2A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \nRST~input (
	.i(nRST),
	.ibar(gnd),
	.o(\nRST~input_o ));
// synopsys translate_off
defparam \nRST~input .bus_hold = "false";
defparam \nRST~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N8
cycloneive_io_ibuf \syif.tbCTRL~input (
	.i(\syif.tbCTRL ),
	.ibar(gnd),
	.o(\syif.tbCTRL~input_o ));
// synopsys translate_off
defparam \syif.tbCTRL~input .bus_hold = "false";
defparam \syif.tbCTRL~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N1
cycloneive_io_ibuf \syif.addr[1]~input (
	.i(\syif.addr [1]),
	.ibar(gnd),
	.o(\syif.addr[1]~input_o ));
// synopsys translate_off
defparam \syif.addr[1]~input .bus_hold = "false";
defparam \syif.addr[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X38_Y73_N15
cycloneive_io_ibuf \syif.addr[0]~input (
	.i(\syif.addr [0]),
	.ibar(gnd),
	.o(\syif.addr[0]~input_o ));
// synopsys translate_off
defparam \syif.addr[0]~input .bus_hold = "false";
defparam \syif.addr[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y44_N15
cycloneive_io_ibuf \syif.addr[3]~input (
	.i(\syif.addr [3]),
	.ibar(gnd),
	.o(\syif.addr[3]~input_o ));
// synopsys translate_off
defparam \syif.addr[3]~input .bus_hold = "false";
defparam \syif.addr[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y42_N1
cycloneive_io_ibuf \syif.addr[2]~input (
	.i(\syif.addr [2]),
	.ibar(gnd),
	.o(\syif.addr[2]~input_o ));
// synopsys translate_off
defparam \syif.addr[2]~input .bus_hold = "false";
defparam \syif.addr[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N22
cycloneive_io_ibuf \syif.addr[5]~input (
	.i(\syif.addr [5]),
	.ibar(gnd),
	.o(\syif.addr[5]~input_o ));
// synopsys translate_off
defparam \syif.addr[5]~input .bus_hold = "false";
defparam \syif.addr[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X38_Y73_N22
cycloneive_io_ibuf \syif.addr[4]~input (
	.i(\syif.addr [4]),
	.ibar(gnd),
	.o(\syif.addr[4]~input_o ));
// synopsys translate_off
defparam \syif.addr[4]~input .bus_hold = "false";
defparam \syif.addr[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X79_Y73_N8
cycloneive_io_ibuf \syif.addr[7]~input (
	.i(\syif.addr [7]),
	.ibar(gnd),
	.o(\syif.addr[7]~input_o ));
// synopsys translate_off
defparam \syif.addr[7]~input .bus_hold = "false";
defparam \syif.addr[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N8
cycloneive_io_ibuf \syif.addr[6]~input (
	.i(\syif.addr [6]),
	.ibar(gnd),
	.o(\syif.addr[6]~input_o ));
// synopsys translate_off
defparam \syif.addr[6]~input .bus_hold = "false";
defparam \syif.addr[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N1
cycloneive_io_ibuf \syif.addr[9]~input (
	.i(\syif.addr [9]),
	.ibar(gnd),
	.o(\syif.addr[9]~input_o ));
// synopsys translate_off
defparam \syif.addr[9]~input .bus_hold = "false";
defparam \syif.addr[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N8
cycloneive_io_ibuf \syif.addr[8]~input (
	.i(\syif.addr [8]),
	.ibar(gnd),
	.o(\syif.addr[8]~input_o ));
// synopsys translate_off
defparam \syif.addr[8]~input .bus_hold = "false";
defparam \syif.addr[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \syif.addr[11]~input (
	.i(\syif.addr [11]),
	.ibar(gnd),
	.o(\syif.addr[11]~input_o ));
// synopsys translate_off
defparam \syif.addr[11]~input .bus_hold = "false";
defparam \syif.addr[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N15
cycloneive_io_ibuf \syif.addr[10]~input (
	.i(\syif.addr [10]),
	.ibar(gnd),
	.o(\syif.addr[10]~input_o ));
// synopsys translate_off
defparam \syif.addr[10]~input .bus_hold = "false";
defparam \syif.addr[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N1
cycloneive_io_ibuf \syif.addr[13]~input (
	.i(\syif.addr [13]),
	.ibar(gnd),
	.o(\syif.addr[13]~input_o ));
// synopsys translate_off
defparam \syif.addr[13]~input .bus_hold = "false";
defparam \syif.addr[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N15
cycloneive_io_ibuf \syif.addr[12]~input (
	.i(\syif.addr [12]),
	.ibar(gnd),
	.o(\syif.addr[12]~input_o ));
// synopsys translate_off
defparam \syif.addr[12]~input .bus_hold = "false";
defparam \syif.addr[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N15
cycloneive_io_ibuf \syif.addr[15]~input (
	.i(\syif.addr [15]),
	.ibar(gnd),
	.o(\syif.addr[15]~input_o ));
// synopsys translate_off
defparam \syif.addr[15]~input .bus_hold = "false";
defparam \syif.addr[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N1
cycloneive_io_ibuf \syif.addr[14]~input (
	.i(\syif.addr [14]),
	.ibar(gnd),
	.o(\syif.addr[14]~input_o ));
// synopsys translate_off
defparam \syif.addr[14]~input .bus_hold = "false";
defparam \syif.addr[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N8
cycloneive_io_ibuf \syif.addr[17]~input (
	.i(\syif.addr [17]),
	.ibar(gnd),
	.o(\syif.addr[17]~input_o ));
// synopsys translate_off
defparam \syif.addr[17]~input .bus_hold = "false";
defparam \syif.addr[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N8
cycloneive_io_ibuf \syif.addr[16]~input (
	.i(\syif.addr [16]),
	.ibar(gnd),
	.o(\syif.addr[16]~input_o ));
// synopsys translate_off
defparam \syif.addr[16]~input .bus_hold = "false";
defparam \syif.addr[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y40_N8
cycloneive_io_ibuf \syif.addr[19]~input (
	.i(\syif.addr [19]),
	.ibar(gnd),
	.o(\syif.addr[19]~input_o ));
// synopsys translate_off
defparam \syif.addr[19]~input .bus_hold = "false";
defparam \syif.addr[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y0_N8
cycloneive_io_ibuf \syif.addr[18]~input (
	.i(\syif.addr [18]),
	.ibar(gnd),
	.o(\syif.addr[18]~input_o ));
// synopsys translate_off
defparam \syif.addr[18]~input .bus_hold = "false";
defparam \syif.addr[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N8
cycloneive_io_ibuf \syif.addr[21]~input (
	.i(\syif.addr [21]),
	.ibar(gnd),
	.o(\syif.addr[21]~input_o ));
// synopsys translate_off
defparam \syif.addr[21]~input .bus_hold = "false";
defparam \syif.addr[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X35_Y73_N22
cycloneive_io_ibuf \syif.addr[20]~input (
	.i(\syif.addr [20]),
	.ibar(gnd),
	.o(\syif.addr[20]~input_o ));
// synopsys translate_off
defparam \syif.addr[20]~input .bus_hold = "false";
defparam \syif.addr[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N15
cycloneive_io_ibuf \syif.addr[23]~input (
	.i(\syif.addr [23]),
	.ibar(gnd),
	.o(\syif.addr[23]~input_o ));
// synopsys translate_off
defparam \syif.addr[23]~input .bus_hold = "false";
defparam \syif.addr[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N15
cycloneive_io_ibuf \syif.addr[22]~input (
	.i(\syif.addr [22]),
	.ibar(gnd),
	.o(\syif.addr[22]~input_o ));
// synopsys translate_off
defparam \syif.addr[22]~input .bus_hold = "false";
defparam \syif.addr[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N15
cycloneive_io_ibuf \syif.addr[25]~input (
	.i(\syif.addr [25]),
	.ibar(gnd),
	.o(\syif.addr[25]~input_o ));
// synopsys translate_off
defparam \syif.addr[25]~input .bus_hold = "false";
defparam \syif.addr[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \syif.addr[24]~input (
	.i(\syif.addr [24]),
	.ibar(gnd),
	.o(\syif.addr[24]~input_o ));
// synopsys translate_off
defparam \syif.addr[24]~input .bus_hold = "false";
defparam \syif.addr[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N8
cycloneive_io_ibuf \syif.addr[27]~input (
	.i(\syif.addr [27]),
	.ibar(gnd),
	.o(\syif.addr[27]~input_o ));
// synopsys translate_off
defparam \syif.addr[27]~input .bus_hold = "false";
defparam \syif.addr[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X38_Y73_N8
cycloneive_io_ibuf \syif.addr[26]~input (
	.i(\syif.addr [26]),
	.ibar(gnd),
	.o(\syif.addr[26]~input_o ));
// synopsys translate_off
defparam \syif.addr[26]~input .bus_hold = "false";
defparam \syif.addr[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N15
cycloneive_io_ibuf \syif.addr[29]~input (
	.i(\syif.addr [29]),
	.ibar(gnd),
	.o(\syif.addr[29]~input_o ));
// synopsys translate_off
defparam \syif.addr[29]~input .bus_hold = "false";
defparam \syif.addr[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N15
cycloneive_io_ibuf \syif.addr[28]~input (
	.i(\syif.addr [28]),
	.ibar(gnd),
	.o(\syif.addr[28]~input_o ));
// synopsys translate_off
defparam \syif.addr[28]~input .bus_hold = "false";
defparam \syif.addr[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N8
cycloneive_io_ibuf \syif.addr[31]~input (
	.i(\syif.addr [31]),
	.ibar(gnd),
	.o(\syif.addr[31]~input_o ));
// synopsys translate_off
defparam \syif.addr[31]~input .bus_hold = "false";
defparam \syif.addr[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N15
cycloneive_io_ibuf \syif.addr[30]~input (
	.i(\syif.addr [30]),
	.ibar(gnd),
	.o(\syif.addr[30]~input_o ));
// synopsys translate_off
defparam \syif.addr[30]~input .bus_hold = "false";
defparam \syif.addr[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N8
cycloneive_io_ibuf \syif.WEN~input (
	.i(\syif.WEN ),
	.ibar(gnd),
	.o(\syif.WEN~input_o ));
// synopsys translate_off
defparam \syif.WEN~input .bus_hold = "false";
defparam \syif.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N8
cycloneive_io_ibuf \syif.REN~input (
	.i(\syif.REN ),
	.ibar(gnd),
	.o(\syif.REN~input_o ));
// synopsys translate_off
defparam \syif.REN~input .bus_hold = "false";
defparam \syif.REN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \CLK~input (
	.i(CLK),
	.ibar(gnd),
	.o(\CLK~input_o ));
// synopsys translate_off
defparam \CLK~input .bus_hold = "false";
defparam \CLK~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y0_N15
cycloneive_io_ibuf \syif.store[0]~input (
	.i(\syif.store [0]),
	.ibar(gnd),
	.o(\syif.store[0]~input_o ));
// synopsys translate_off
defparam \syif.store[0]~input .bus_hold = "false";
defparam \syif.store[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N22
cycloneive_io_ibuf \syif.store[1]~input (
	.i(\syif.store [1]),
	.ibar(gnd),
	.o(\syif.store[1]~input_o ));
// synopsys translate_off
defparam \syif.store[1]~input .bus_hold = "false";
defparam \syif.store[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N1
cycloneive_io_ibuf \syif.store[2]~input (
	.i(\syif.store [2]),
	.ibar(gnd),
	.o(\syif.store[2]~input_o ));
// synopsys translate_off
defparam \syif.store[2]~input .bus_hold = "false";
defparam \syif.store[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y0_N22
cycloneive_io_ibuf \syif.store[3]~input (
	.i(\syif.store [3]),
	.ibar(gnd),
	.o(\syif.store[3]~input_o ));
// synopsys translate_off
defparam \syif.store[3]~input .bus_hold = "false";
defparam \syif.store[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N1
cycloneive_io_ibuf \syif.store[4]~input (
	.i(\syif.store [4]),
	.ibar(gnd),
	.o(\syif.store[4]~input_o ));
// synopsys translate_off
defparam \syif.store[4]~input .bus_hold = "false";
defparam \syif.store[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N22
cycloneive_io_ibuf \syif.store[5]~input (
	.i(\syif.store [5]),
	.ibar(gnd),
	.o(\syif.store[5]~input_o ));
// synopsys translate_off
defparam \syif.store[5]~input .bus_hold = "false";
defparam \syif.store[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N15
cycloneive_io_ibuf \syif.store[6]~input (
	.i(\syif.store [6]),
	.ibar(gnd),
	.o(\syif.store[6]~input_o ));
// synopsys translate_off
defparam \syif.store[6]~input .bus_hold = "false";
defparam \syif.store[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N22
cycloneive_io_ibuf \syif.store[7]~input (
	.i(\syif.store [7]),
	.ibar(gnd),
	.o(\syif.store[7]~input_o ));
// synopsys translate_off
defparam \syif.store[7]~input .bus_hold = "false";
defparam \syif.store[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N1
cycloneive_io_ibuf \syif.store[8]~input (
	.i(\syif.store [8]),
	.ibar(gnd),
	.o(\syif.store[8]~input_o ));
// synopsys translate_off
defparam \syif.store[8]~input .bus_hold = "false";
defparam \syif.store[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N8
cycloneive_io_ibuf \syif.store[9]~input (
	.i(\syif.store [9]),
	.ibar(gnd),
	.o(\syif.store[9]~input_o ));
// synopsys translate_off
defparam \syif.store[9]~input .bus_hold = "false";
defparam \syif.store[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y42_N15
cycloneive_io_ibuf \syif.store[10]~input (
	.i(\syif.store [10]),
	.ibar(gnd),
	.o(\syif.store[10]~input_o ));
// synopsys translate_off
defparam \syif.store[10]~input .bus_hold = "false";
defparam \syif.store[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N1
cycloneive_io_ibuf \syif.store[11]~input (
	.i(\syif.store [11]),
	.ibar(gnd),
	.o(\syif.store[11]~input_o ));
// synopsys translate_off
defparam \syif.store[11]~input .bus_hold = "false";
defparam \syif.store[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N8
cycloneive_io_ibuf \syif.store[12]~input (
	.i(\syif.store [12]),
	.ibar(gnd),
	.o(\syif.store[12]~input_o ));
// synopsys translate_off
defparam \syif.store[12]~input .bus_hold = "false";
defparam \syif.store[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N15
cycloneive_io_ibuf \syif.store[13]~input (
	.i(\syif.store [13]),
	.ibar(gnd),
	.o(\syif.store[13]~input_o ));
// synopsys translate_off
defparam \syif.store[13]~input .bus_hold = "false";
defparam \syif.store[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N1
cycloneive_io_ibuf \syif.store[14]~input (
	.i(\syif.store [14]),
	.ibar(gnd),
	.o(\syif.store[14]~input_o ));
// synopsys translate_off
defparam \syif.store[14]~input .bus_hold = "false";
defparam \syif.store[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N22
cycloneive_io_ibuf \syif.store[15]~input (
	.i(\syif.store [15]),
	.ibar(gnd),
	.o(\syif.store[15]~input_o ));
// synopsys translate_off
defparam \syif.store[15]~input .bus_hold = "false";
defparam \syif.store[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N15
cycloneive_io_ibuf \syif.store[16]~input (
	.i(\syif.store [16]),
	.ibar(gnd),
	.o(\syif.store[16]~input_o ));
// synopsys translate_off
defparam \syif.store[16]~input .bus_hold = "false";
defparam \syif.store[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N22
cycloneive_io_ibuf \syif.store[17]~input (
	.i(\syif.store [17]),
	.ibar(gnd),
	.o(\syif.store[17]~input_o ));
// synopsys translate_off
defparam \syif.store[17]~input .bus_hold = "false";
defparam \syif.store[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y73_N22
cycloneive_io_ibuf \syif.store[18]~input (
	.i(\syif.store [18]),
	.ibar(gnd),
	.o(\syif.store[18]~input_o ));
// synopsys translate_off
defparam \syif.store[18]~input .bus_hold = "false";
defparam \syif.store[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N22
cycloneive_io_ibuf \syif.store[19]~input (
	.i(\syif.store [19]),
	.ibar(gnd),
	.o(\syif.store[19]~input_o ));
// synopsys translate_off
defparam \syif.store[19]~input .bus_hold = "false";
defparam \syif.store[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N15
cycloneive_io_ibuf \syif.store[20]~input (
	.i(\syif.store [20]),
	.ibar(gnd),
	.o(\syif.store[20]~input_o ));
// synopsys translate_off
defparam \syif.store[20]~input .bus_hold = "false";
defparam \syif.store[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N8
cycloneive_io_ibuf \syif.store[21]~input (
	.i(\syif.store [21]),
	.ibar(gnd),
	.o(\syif.store[21]~input_o ));
// synopsys translate_off
defparam \syif.store[21]~input .bus_hold = "false";
defparam \syif.store[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N1
cycloneive_io_ibuf \syif.store[22]~input (
	.i(\syif.store [22]),
	.ibar(gnd),
	.o(\syif.store[22]~input_o ));
// synopsys translate_off
defparam \syif.store[22]~input .bus_hold = "false";
defparam \syif.store[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N22
cycloneive_io_ibuf \syif.store[23]~input (
	.i(\syif.store [23]),
	.ibar(gnd),
	.o(\syif.store[23]~input_o ));
// synopsys translate_off
defparam \syif.store[23]~input .bus_hold = "false";
defparam \syif.store[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N1
cycloneive_io_ibuf \syif.store[24]~input (
	.i(\syif.store [24]),
	.ibar(gnd),
	.o(\syif.store[24]~input_o ));
// synopsys translate_off
defparam \syif.store[24]~input .bus_hold = "false";
defparam \syif.store[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N22
cycloneive_io_ibuf \syif.store[25]~input (
	.i(\syif.store [25]),
	.ibar(gnd),
	.o(\syif.store[25]~input_o ));
// synopsys translate_off
defparam \syif.store[25]~input .bus_hold = "false";
defparam \syif.store[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N15
cycloneive_io_ibuf \syif.store[26]~input (
	.i(\syif.store [26]),
	.ibar(gnd),
	.o(\syif.store[26]~input_o ));
// synopsys translate_off
defparam \syif.store[26]~input .bus_hold = "false";
defparam \syif.store[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N22
cycloneive_io_ibuf \syif.store[27]~input (
	.i(\syif.store [27]),
	.ibar(gnd),
	.o(\syif.store[27]~input_o ));
// synopsys translate_off
defparam \syif.store[27]~input .bus_hold = "false";
defparam \syif.store[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N1
cycloneive_io_ibuf \syif.store[28]~input (
	.i(\syif.store [28]),
	.ibar(gnd),
	.o(\syif.store[28]~input_o ));
// synopsys translate_off
defparam \syif.store[28]~input .bus_hold = "false";
defparam \syif.store[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y41_N8
cycloneive_io_ibuf \syif.store[29]~input (
	.i(\syif.store [29]),
	.ibar(gnd),
	.o(\syif.store[29]~input_o ));
// synopsys translate_off
defparam \syif.store[29]~input .bus_hold = "false";
defparam \syif.store[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N1
cycloneive_io_ibuf \syif.store[30]~input (
	.i(\syif.store [30]),
	.ibar(gnd),
	.o(\syif.store[30]~input_o ));
// synopsys translate_off
defparam \syif.store[30]~input .bus_hold = "false";
defparam \syif.store[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y40_N1
cycloneive_io_ibuf \syif.store[31]~input (
	.i(\syif.store [31]),
	.ibar(gnd),
	.o(\syif.store[31]~input_o ));
// synopsys translate_off
defparam \syif.store[31]~input .bus_hold = "false";
defparam \syif.store[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G4
cycloneive_clkctrl \altera_internal_jtag~TCKUTAPclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\altera_internal_jtag~TCKUTAP }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
// synopsys translate_off
defparam \altera_internal_jtag~TCKUTAPclkctrl .clock_type = "global clock";
defparam \altera_internal_jtag~TCKUTAPclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G7
cycloneive_clkctrl \CPUCLK~clkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CPUCLK~q }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CPUCLK~clkctrl_outclk ));
// synopsys translate_off
defparam \CPUCLK~clkctrl .clock_type = "global clock";
defparam \CPUCLK~clkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G1
cycloneive_clkctrl \nRST~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\nRST~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\nRST~inputclkctrl_outclk ));
// synopsys translate_off
defparam \nRST~inputclkctrl .clock_type = "global clock";
defparam \nRST~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \CLK~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CLK~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CLK~inputclkctrl_outclk ));
// synopsys translate_off
defparam \CLK~inputclkctrl .clock_type = "global clock";
defparam \CLK~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOOBUF_X0_Y31_N16
cycloneive_io_obuf \syif.halt~output (
	.i(\CPU|DP|dpif.halt~q ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.halt ),
	.obar());
// synopsys translate_off
defparam \syif.halt~output .bus_hold = "false";
defparam \syif.halt~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N9
cycloneive_io_obuf \syif.load[0]~output (
	.i(\RAM|ramif.ramload[0]~1_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [0]),
	.obar());
// synopsys translate_off
defparam \syif.load[0]~output .bus_hold = "false";
defparam \syif.load[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N2
cycloneive_io_obuf \syif.load[1]~output (
	.i(\RAM|ramif.ramload[1]~2_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [1]),
	.obar());
// synopsys translate_off
defparam \syif.load[1]~output .bus_hold = "false";
defparam \syif.load[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N2
cycloneive_io_obuf \syif.load[2]~output (
	.i(\RAM|ramif.ramload[2]~4_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [2]),
	.obar());
// synopsys translate_off
defparam \syif.load[2]~output .bus_hold = "false";
defparam \syif.load[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X72_Y73_N23
cycloneive_io_obuf \syif.load[3]~output (
	.i(\RAM|ramif.ramload[3]~5_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [3]),
	.obar());
// synopsys translate_off
defparam \syif.load[3]~output .bus_hold = "false";
defparam \syif.load[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N2
cycloneive_io_obuf \syif.load[4]~output (
	.i(\RAM|ramif.ramload[4]~7_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [4]),
	.obar());
// synopsys translate_off
defparam \syif.load[4]~output .bus_hold = "false";
defparam \syif.load[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X69_Y73_N16
cycloneive_io_obuf \syif.load[5]~output (
	.i(\RAM|ramif.ramload[5]~9_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [5]),
	.obar());
// synopsys translate_off
defparam \syif.load[5]~output .bus_hold = "false";
defparam \syif.load[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N23
cycloneive_io_obuf \syif.load[6]~output (
	.i(\RAM|ramif.ramload[6]~10_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [6]),
	.obar());
// synopsys translate_off
defparam \syif.load[6]~output .bus_hold = "false";
defparam \syif.load[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N23
cycloneive_io_obuf \syif.load[7]~output (
	.i(\RAM|ramif.ramload[7]~11_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [7]),
	.obar());
// synopsys translate_off
defparam \syif.load[7]~output .bus_hold = "false";
defparam \syif.load[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N2
cycloneive_io_obuf \syif.load[8]~output (
	.i(\RAM|ramif.ramload[8]~12_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [8]),
	.obar());
// synopsys translate_off
defparam \syif.load[8]~output .bus_hold = "false";
defparam \syif.load[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N16
cycloneive_io_obuf \syif.load[9]~output (
	.i(\RAM|ramif.ramload[9]~13_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [9]),
	.obar());
// synopsys translate_off
defparam \syif.load[9]~output .bus_hold = "false";
defparam \syif.load[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X74_Y73_N16
cycloneive_io_obuf \syif.load[10]~output (
	.i(\RAM|ramif.ramload[10]~14_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [10]),
	.obar());
// synopsys translate_off
defparam \syif.load[10]~output .bus_hold = "false";
defparam \syif.load[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N9
cycloneive_io_obuf \syif.load[11]~output (
	.i(\RAM|ramif.ramload[11]~15_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [11]),
	.obar());
// synopsys translate_off
defparam \syif.load[11]~output .bus_hold = "false";
defparam \syif.load[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y73_N16
cycloneive_io_obuf \syif.load[12]~output (
	.i(\RAM|ramif.ramload[12]~16_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [12]),
	.obar());
// synopsys translate_off
defparam \syif.load[12]~output .bus_hold = "false";
defparam \syif.load[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N2
cycloneive_io_obuf \syif.load[13]~output (
	.i(\RAM|ramif.ramload[13]~17_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [13]),
	.obar());
// synopsys translate_off
defparam \syif.load[13]~output .bus_hold = "false";
defparam \syif.load[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N9
cycloneive_io_obuf \syif.load[14]~output (
	.i(\RAM|ramif.ramload[14]~18_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [14]),
	.obar());
// synopsys translate_off
defparam \syif.load[14]~output .bus_hold = "false";
defparam \syif.load[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N9
cycloneive_io_obuf \syif.load[15]~output (
	.i(\RAM|ramif.ramload[15]~19_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [15]),
	.obar());
// synopsys translate_off
defparam \syif.load[15]~output .bus_hold = "false";
defparam \syif.load[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y35_N2
cycloneive_io_obuf \syif.load[16]~output (
	.i(\RAM|ramif.ramload[16]~21_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [16]),
	.obar());
// synopsys translate_off
defparam \syif.load[16]~output .bus_hold = "false";
defparam \syif.load[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y34_N2
cycloneive_io_obuf \syif.load[17]~output (
	.i(\RAM|ramif.ramload[17]~23_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [17]),
	.obar());
// synopsys translate_off
defparam \syif.load[17]~output .bus_hold = "false";
defparam \syif.load[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y73_N2
cycloneive_io_obuf \syif.load[18]~output (
	.i(\RAM|ramif.ramload[18]~24_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [18]),
	.obar());
// synopsys translate_off
defparam \syif.load[18]~output .bus_hold = "false";
defparam \syif.load[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y73_N23
cycloneive_io_obuf \syif.load[19]~output (
	.i(\RAM|ramif.ramload[19]~25_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [19]),
	.obar());
// synopsys translate_off
defparam \syif.load[19]~output .bus_hold = "false";
defparam \syif.load[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X45_Y0_N16
cycloneive_io_obuf \syif.load[20]~output (
	.i(\RAM|ramif.ramload[20]~26_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [20]),
	.obar());
// synopsys translate_off
defparam \syif.load[20]~output .bus_hold = "false";
defparam \syif.load[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X42_Y73_N2
cycloneive_io_obuf \syif.load[21]~output (
	.i(\RAM|ramif.ramload[21]~27_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [21]),
	.obar());
// synopsys translate_off
defparam \syif.load[21]~output .bus_hold = "false";
defparam \syif.load[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y43_N16
cycloneive_io_obuf \syif.load[22]~output (
	.i(\RAM|ramif.ramload[22]~28_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [22]),
	.obar());
// synopsys translate_off
defparam \syif.load[22]~output .bus_hold = "false";
defparam \syif.load[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N16
cycloneive_io_obuf \syif.load[23]~output (
	.i(\RAM|ramif.ramload[23]~29_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [23]),
	.obar());
// synopsys translate_off
defparam \syif.load[23]~output .bus_hold = "false";
defparam \syif.load[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y0_N2
cycloneive_io_obuf \syif.load[24]~output (
	.i(\RAM|ramif.ramload[24]~30_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [24]),
	.obar());
// synopsys translate_off
defparam \syif.load[24]~output .bus_hold = "false";
defparam \syif.load[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N9
cycloneive_io_obuf \syif.load[25]~output (
	.i(\RAM|ramif.ramload[25]~31_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [25]),
	.obar());
// synopsys translate_off
defparam \syif.load[25]~output .bus_hold = "false";
defparam \syif.load[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N9
cycloneive_io_obuf \syif.load[26]~output (
	.i(\RAM|ramif.ramload[26]~33_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [26]),
	.obar());
// synopsys translate_off
defparam \syif.load[26]~output .bus_hold = "false";
defparam \syif.load[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X72_Y73_N16
cycloneive_io_obuf \syif.load[27]~output (
	.i(\RAM|ramif.ramload[27]~35_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [27]),
	.obar());
// synopsys translate_off
defparam \syif.load[27]~output .bus_hold = "false";
defparam \syif.load[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N16
cycloneive_io_obuf \syif.load[28]~output (
	.i(\RAM|ramif.ramload[28]~37_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [28]),
	.obar());
// synopsys translate_off
defparam \syif.load[28]~output .bus_hold = "false";
defparam \syif.load[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y42_N9
cycloneive_io_obuf \syif.load[29]~output (
	.i(\RAM|ramif.ramload[29]~39_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [29]),
	.obar());
// synopsys translate_off
defparam \syif.load[29]~output .bus_hold = "false";
defparam \syif.load[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N9
cycloneive_io_obuf \syif.load[30]~output (
	.i(\RAM|ramif.ramload[30]~41_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [30]),
	.obar());
// synopsys translate_off
defparam \syif.load[30]~output .bus_hold = "false";
defparam \syif.load[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y73_N2
cycloneive_io_obuf \syif.load[31]~output (
	.i(\RAM|ramif.ramload[31]~43_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [31]),
	.obar());
// synopsys translate_off
defparam \syif.load[31]~output .bus_hold = "false";
defparam \syif.load[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y37_N1
cycloneive_io_obuf \altera_reserved_tdo~output (
	.i(\altera_internal_jtag~TDO ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(altera_reserved_tdo),
	.obar());
// synopsys translate_off
defparam \altera_reserved_tdo~output .bus_hold = "false";
defparam \altera_reserved_tdo~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y38_N1
cycloneive_io_ibuf \altera_reserved_tms~input (
	.i(altera_reserved_tms),
	.ibar(gnd),
	.o(\altera_reserved_tms~input_o ));
// synopsys translate_off
defparam \altera_reserved_tms~input .bus_hold = "false";
defparam \altera_reserved_tms~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y39_N1
cycloneive_io_ibuf \altera_reserved_tck~input (
	.i(altera_reserved_tck),
	.ibar(gnd),
	.o(\altera_reserved_tck~input_o ));
// synopsys translate_off
defparam \altera_reserved_tck~input .bus_hold = "false";
defparam \altera_reserved_tck~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y40_N1
cycloneive_io_ibuf \altera_reserved_tdi~input (
	.i(altera_reserved_tdi),
	.ibar(gnd),
	.o(\altera_reserved_tdi~input_o ));
// synopsys translate_off
defparam \altera_reserved_tdi~input .bus_hold = "false";
defparam \altera_reserved_tdi~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .lut_mask = 16'hE0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .lut_mask = 16'hFFFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .lut_mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N22
cycloneive_lcell_comb \~QIC_CREATED_GND~I (
// Equation(s):
// \~QIC_CREATED_GND~I_combout  = GND

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
// synopsys translate_off
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y39_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .lut_mask = 16'h3373;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y39_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y39_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .lut_mask = 16'hFFFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y39_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .lut_mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .lut_mask = 16'h1000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .lut_mask = 16'hA080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .lut_mask = 16'h22F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .lut_mask = 16'hF0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .lut_mask = 16'hFFFB;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y39_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .lut_mask = 16'hAAA8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .lut_mask = 16'hFA0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .lut_mask = 16'hFA50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .lut_mask = 16'h00A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .lut_mask = 16'h7250;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .lut_mask = 16'hCFC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .lut_mask = 16'hEE44;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .lut_mask = 16'hC808;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .lut_mask = 16'hE4E4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .lut_mask = 16'hFC0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .lut_mask = 16'hFC0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .lut_mask = 16'hFC0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .lut_mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .lut_mask = 16'hFC22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .lut_mask = 16'hD9C8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .lut_mask = 16'hC8D8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .lut_mask = 16'hFAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .lut_mask = 16'h07F3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y36_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.clk(!\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X12_Y38_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X17_Y4_N0
cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ram (
	is_in_use_reg,
	ramiframload_0,
	LessThan1,
	ramaddr,
	ramaddr1,
	ramaddr2,
	ramaddr3,
	ramaddr4,
	ramaddr5,
	ramaddr6,
	ramaddr7,
	always0,
	ramaddr8,
	ramaddr9,
	ramaddr10,
	ramaddr11,
	ramaddr12,
	ramaddr13,
	ramaddr14,
	ramaddr15,
	always01,
	ramaddr16,
	ramaddr17,
	\ramif.ramaddr ,
	ramaddr18,
	ramaddr19,
	ramaddr20,
	ramaddr21,
	ramaddr22,
	ramaddr23,
	ramaddr24,
	ramaddr25,
	ramaddr26,
	ramaddr27,
	ramaddr28,
	ramaddr29,
	\ramif.ramWEN ,
	\ramif.ramREN ,
	always02,
	always03,
	ramiframload_01,
	always1,
	ramiframload_1,
	ramiframload_2,
	ramiframload_21,
	ramiframload_3,
	ramiframload_4,
	ramiframload_41,
	ramiframload_5,
	ramiframload_51,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_161,
	ramiframload_17,
	ramiframload_171,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_211,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_261,
	ramiframload_27,
	ramiframload_271,
	ramiframload_28,
	ramiframload_281,
	ramiframload_29,
	ramiframload_291,
	ramiframload_30,
	ramiframload_301,
	ramiframload_31,
	ramiframload_311,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramstore,
	ramstore1,
	ramstore2,
	ramstore3,
	ramstore4,
	ramstore5,
	ramstore6,
	ramstore7,
	ramstore8,
	ramstore9,
	ramstore10,
	ramstore11,
	ramstore12,
	ramstore13,
	ramstore14,
	ramstore15,
	ramstore16,
	ramstore17,
	ramstore18,
	ramstore19,
	ramstore20,
	ramstore21,
	ramstore22,
	ramstore23,
	ramstore24,
	ramstore25,
	ramstore26,
	ramstore27,
	ramstore28,
	ramstore29,
	ramstore30,
	ramstore31,
	ramaddr30,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	nRST,
	altera_internal_jtag1,
	nRST1,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	is_in_use_reg;
output 	ramiframload_0;
output 	LessThan1;
input 	ramaddr;
input 	ramaddr1;
input 	ramaddr2;
input 	ramaddr3;
input 	ramaddr4;
input 	ramaddr5;
input 	ramaddr6;
input 	ramaddr7;
output 	always0;
input 	ramaddr8;
input 	ramaddr9;
input 	ramaddr10;
input 	ramaddr11;
input 	ramaddr12;
input 	ramaddr13;
input 	ramaddr14;
input 	ramaddr15;
output 	always01;
input 	ramaddr16;
input 	ramaddr17;
input 	[31:0] \ramif.ramaddr ;
input 	ramaddr18;
input 	ramaddr19;
input 	ramaddr20;
input 	ramaddr21;
input 	ramaddr22;
input 	ramaddr23;
input 	ramaddr24;
input 	ramaddr25;
input 	ramaddr26;
input 	ramaddr27;
input 	ramaddr28;
input 	ramaddr29;
input 	\ramif.ramWEN ;
input 	\ramif.ramREN ;
output 	always02;
output 	always03;
output 	ramiframload_01;
output 	always1;
output 	ramiframload_1;
output 	ramiframload_2;
output 	ramiframload_21;
output 	ramiframload_3;
output 	ramiframload_4;
output 	ramiframload_41;
output 	ramiframload_5;
output 	ramiframload_51;
output 	ramiframload_6;
output 	ramiframload_7;
output 	ramiframload_8;
output 	ramiframload_9;
output 	ramiframload_10;
output 	ramiframload_11;
output 	ramiframload_12;
output 	ramiframload_13;
output 	ramiframload_14;
output 	ramiframload_15;
output 	ramiframload_16;
output 	ramiframload_161;
output 	ramiframload_17;
output 	ramiframload_171;
output 	ramiframload_18;
output 	ramiframload_19;
output 	ramiframload_20;
output 	ramiframload_211;
output 	ramiframload_22;
output 	ramiframload_23;
output 	ramiframload_24;
output 	ramiframload_25;
output 	ramiframload_26;
output 	ramiframload_261;
output 	ramiframload_27;
output 	ramiframload_271;
output 	ramiframload_28;
output 	ramiframload_281;
output 	ramiframload_29;
output 	ramiframload_291;
output 	ramiframload_30;
output 	ramiframload_301;
output 	ramiframload_31;
output 	ramiframload_311;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramstore;
input 	ramstore1;
input 	ramstore2;
input 	ramstore3;
input 	ramstore4;
input 	ramstore5;
input 	ramstore6;
input 	ramstore7;
input 	ramstore8;
input 	ramstore9;
input 	ramstore10;
input 	ramstore11;
input 	ramstore12;
input 	ramstore13;
input 	ramstore14;
input 	ramstore15;
input 	ramstore16;
input 	ramstore17;
input 	ramstore18;
input 	ramstore19;
input 	ramstore20;
input 	ramstore21;
input 	ramstore22;
input 	ramstore23;
input 	ramstore24;
input 	ramstore25;
input 	ramstore26;
input 	ramstore27;
input 	ramstore28;
input 	ramstore29;
input 	ramstore30;
input 	ramstore31;
input 	ramaddr30;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	nRST;
input 	altera_internal_jtag1;
input 	nRST1;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ;
wire \addr[21]~feeder_combout ;
wire \addr[23]~feeder_combout ;
wire \addr[27]~feeder_combout ;
wire \addr[29]~feeder_combout ;
wire \always0~22_combout ;
wire \always0~23_combout ;
wire \count[1]~2_combout ;
wire \LessThan1~1_combout ;
wire \count[2]~1_combout ;
wire \count[0]~3_combout ;
wire \count[3]~0_combout ;
wire \always0~1_combout ;
wire \always0~0_combout ;
wire \addr[5]~feeder_combout ;
wire \always0~2_combout ;
wire \addr[7]~feeder_combout ;
wire \always0~3_combout ;
wire \always0~5_combout ;
wire \always0~8_combout ;
wire \addr[11]~feeder_combout ;
wire \always0~6_combout ;
wire \addr[13]~feeder_combout ;
wire \always0~7_combout ;
wire \always0~16_combout ;
wire \always0~18_combout ;
wire \addr[25]~feeder_combout ;
wire \always0~15_combout ;
wire \always0~17_combout ;
wire \always0~19_combout ;
wire \always0~11_combout ;
wire \always0~12_combout ;
wire \always0~10_combout ;
wire \always0~13_combout ;
wire \always0~14_combout ;
wire \always1~0_combout ;
wire [1:0] en;
wire [3:0] count;
wire [31:0] addr;
wire [0:0] \altsyncram_component|auto_generated|altsyncram1|address_reg_a ;


altsyncram_1 altsyncram_component(
	.ram_block3a32(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.ram_block3a0(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.ram_block3a33(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.ram_block3a1(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.ram_block3a34(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.ram_block3a2(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.ram_block3a35(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.ram_block3a3(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.ram_block3a36(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.ram_block3a4(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.ram_block3a37(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.ram_block3a5(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.ram_block3a38(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.ram_block3a6(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.ram_block3a39(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.ram_block3a7(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.ram_block3a40(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.ram_block3a8(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.ram_block3a41(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.ram_block3a9(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.ram_block3a42(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.ram_block3a10(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.ram_block3a43(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.ram_block3a11(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.ram_block3a44(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.ram_block3a12(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.ram_block3a45(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.ram_block3a13(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.ram_block3a46(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.ram_block3a14(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.ram_block3a47(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.ram_block3a15(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.ram_block3a48(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.ram_block3a16(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.ram_block3a49(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.ram_block3a17(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.ram_block3a50(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.ram_block3a18(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.ram_block3a51(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.ram_block3a19(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.ram_block3a52(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.ram_block3a20(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.ram_block3a53(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.ram_block3a21(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.ram_block3a54(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.ram_block3a22(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.ram_block3a55(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.ram_block3a23(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.ram_block3a56(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.ram_block3a24(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.ram_block3a57(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.ram_block3a25(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.ram_block3a58(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.ram_block3a26(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.ram_block3a59(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.ram_block3a27(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.ram_block3a60(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.ram_block3a28(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.ram_block3a61(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.ram_block3a29(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.ram_block3a62(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.ram_block3a30(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.ram_block3a63(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.ram_block3a31(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.address_a({gnd,ramaddr15,ramaddr12,ramaddr13,ramaddr10,ramaddr11,ramaddr8,ramaddr9,ramaddr6,ramaddr7,ramaddr4,ramaddr5,ramaddr2,ramaddr3}),
	.ramaddr(ramaddr14),
	.ramWEN(\ramif.ramWEN ),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({ramstore31,ramstore30,ramstore29,ramstore28,ramstore27,ramstore26,ramstore25,ramstore24,ramstore23,ramstore22,ramstore21,ramstore20,ramstore19,ramstore18,ramstore17,ramstore16,ramstore15,ramstore14,ramstore13,ramstore12,ramstore11,ramstore10,ramstore9,ramstore8,ramstore7,ramstore6,
ramstore5,ramstore4,ramstore3,ramstore2,ramstore1,ramstore}),
	.ramaddr1(ramaddr30),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X56_Y39_N23
dffeas \addr[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr16),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[17] .is_wysiwyg = "true";
defparam \addr[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N23
dffeas \addr[21] (
	.clk(CLK),
	.d(\addr[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[21] .is_wysiwyg = "true";
defparam \addr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y43_N15
dffeas \addr[23] (
	.clk(CLK),
	.d(\addr[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[23] .is_wysiwyg = "true";
defparam \addr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N29
dffeas \addr[27] (
	.clk(CLK),
	.d(\addr[27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[27] .is_wysiwyg = "true";
defparam \addr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N23
dffeas \addr[29] (
	.clk(CLK),
	.d(\addr[29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[29] .is_wysiwyg = "true";
defparam \addr[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N22
cycloneive_lcell_comb \addr[21]~feeder (
// Equation(s):
// \addr[21]~feeder_combout  = \ramaddr~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr19),
	.cin(gnd),
	.combout(\addr[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[21]~feeder .lut_mask = 16'hFF00;
defparam \addr[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N14
cycloneive_lcell_comb \addr[23]~feeder (
// Equation(s):
// \addr[23]~feeder_combout  = \ramaddr~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr21),
	.cin(gnd),
	.combout(\addr[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[23]~feeder .lut_mask = 16'hFF00;
defparam \addr[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N28
cycloneive_lcell_comb \addr[27]~feeder (
// Equation(s):
// \addr[27]~feeder_combout  = \ramaddr~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr25),
	.cin(gnd),
	.combout(\addr[27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[27]~feeder .lut_mask = 16'hFF00;
defparam \addr[27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N22
cycloneive_lcell_comb \addr[29]~feeder (
// Equation(s):
// \addr[29]~feeder_combout  = \ramaddr~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr27),
	.cin(gnd),
	.combout(\addr[29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[29]~feeder .lut_mask = 16'hFF00;
defparam \addr[29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N20
cycloneive_lcell_comb \ramif.ramload[0]~0 (
// Equation(s):
// ramiframload_0 = (address_reg_a_0 & (ram_block3a321)) # (!address_reg_a_0 & ((ram_block3a01)))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(gnd),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.cin(gnd),
	.combout(ramiframload_0),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~0 .lut_mask = 16'hF5A0;
defparam \ramif.ramload[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N8
cycloneive_lcell_comb \LessThan1~0 (
// Equation(s):
// LessThan1 = (count[2]) # ((count[3]) # ((count[1] & count[0])))

	.dataa(count[1]),
	.datab(count[2]),
	.datac(count[0]),
	.datad(count[3]),
	.cin(gnd),
	.combout(LessThan1),
	.cout());
// synopsys translate_off
defparam \LessThan1~0 .lut_mask = 16'hFFEC;
defparam \LessThan1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N26
cycloneive_lcell_comb \always0~4 (
// Equation(s):
// always0 = (\always0~1_combout  & (\always0~0_combout  & (\always0~2_combout  & \always0~3_combout )))

	.dataa(\always0~1_combout ),
	.datab(\always0~0_combout ),
	.datac(\always0~2_combout ),
	.datad(\always0~3_combout ),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~4 .lut_mask = 16'h8000;
defparam \always0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N20
cycloneive_lcell_comb \always0~9 (
// Equation(s):
// always01 = (\always0~5_combout  & (\always0~8_combout  & (\always0~6_combout  & \always0~7_combout )))

	.dataa(\always0~5_combout ),
	.datab(\always0~8_combout ),
	.datac(\always0~6_combout ),
	.datad(\always0~7_combout ),
	.cin(gnd),
	.combout(always01),
	.cout());
// synopsys translate_off
defparam \always0~9 .lut_mask = 16'h8000;
defparam \always0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N30
cycloneive_lcell_comb \always0~20 (
// Equation(s):
// always02 = (\always0~19_combout  & (\always0~14_combout  & ((!\ramWEN~0_combout ) # (!\ramREN~1_combout ))))

	.dataa(\ramif.ramREN ),
	.datab(\ramif.ramWEN ),
	.datac(\always0~19_combout ),
	.datad(\always0~14_combout ),
	.cin(gnd),
	.combout(always02),
	.cout());
// synopsys translate_off
defparam \always0~20 .lut_mask = 16'h7000;
defparam \always0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N28
cycloneive_lcell_comb \always0~21 (
// Equation(s):
// always03 = (always0 & (always02 & always01))

	.dataa(always0),
	.datab(always02),
	.datac(gnd),
	.datad(always01),
	.cin(gnd),
	.combout(always03),
	.cout());
// synopsys translate_off
defparam \always0~21 .lut_mask = 16'h8800;
defparam \always0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N20
cycloneive_lcell_comb \ramif.ramload[0]~1 (
// Equation(s):
// ramiframload_01 = (ramiframload_0) # ((\nRST~input_o  & ((!LessThan1) # (!always03))))

	.dataa(ramiframload_0),
	.datab(always03),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(ramiframload_01),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~1 .lut_mask = 16'hBFAA;
defparam \ramif.ramload[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N22
cycloneive_lcell_comb \always1~1 (
// Equation(s):
// always1 = ((always0 & (always02 & \always1~0_combout ))) # (!\nRST~input_o )

	.dataa(always0),
	.datab(nRST),
	.datac(always02),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~1 .lut_mask = 16'hB333;
defparam \always1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N8
cycloneive_lcell_comb \ramif.ramload[1]~2 (
// Equation(s):
// ramiframload_1 = (always1 & ((address_reg_a_0 & (ram_block3a331)) # (!address_reg_a_0 & ((ram_block3a110)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_1),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~2 .lut_mask = 16'hB800;
defparam \ramif.ramload[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N6
cycloneive_lcell_comb \ramif.ramload[2]~3 (
// Equation(s):
// ramiframload_2 = (address_reg_a_0 & ((ram_block3a341))) # (!address_reg_a_0 & (ram_block3a210))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(gnd),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.cin(gnd),
	.combout(ramiframload_2),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~3 .lut_mask = 16'hEE22;
defparam \ramif.ramload[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N14
cycloneive_lcell_comb \ramif.ramload[2]~4 (
// Equation(s):
// ramiframload_21 = (ramiframload_2 & (((LessThan1 & always03)) # (!\nRST~input_o )))

	.dataa(ramiframload_2),
	.datab(nRST),
	.datac(LessThan1),
	.datad(always03),
	.cin(gnd),
	.combout(ramiframload_21),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~4 .lut_mask = 16'hA222;
defparam \ramif.ramload[2]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N24
cycloneive_lcell_comb \ramif.ramload[3]~5 (
// Equation(s):
// ramiframload_3 = (always1 & ((address_reg_a_0 & (ram_block3a351)) # (!address_reg_a_0 & ((ram_block3a310)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.cin(gnd),
	.combout(ramiframload_3),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[3]~5 .lut_mask = 16'hA280;
defparam \ramif.ramload[3]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N18
cycloneive_lcell_comb \ramif.ramload[4]~6 (
// Equation(s):
// ramiframload_4 = (address_reg_a_0 & ((ram_block3a361))) # (!address_reg_a_0 & (ram_block3a410))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.cin(gnd),
	.combout(ramiframload_4),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~6 .lut_mask = 16'hFC30;
defparam \ramif.ramload[4]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N4
cycloneive_lcell_comb \ramif.ramload[4]~7 (
// Equation(s):
// ramiframload_41 = (ramiframload_4) # ((\nRST~input_o  & ((!LessThan1) # (!always03))))

	.dataa(always03),
	.datab(ramiframload_4),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(ramiframload_41),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~7 .lut_mask = 16'hDFCC;
defparam \ramif.ramload[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N16
cycloneive_lcell_comb \ramif.ramload[5]~8 (
// Equation(s):
// ramiframload_5 = (address_reg_a_0 & ((ram_block3a371))) # (!address_reg_a_0 & (ram_block3a510))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(gnd),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.cin(gnd),
	.combout(ramiframload_5),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~8 .lut_mask = 16'hFA50;
defparam \ramif.ramload[5]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N10
cycloneive_lcell_comb \ramif.ramload[5]~9 (
// Equation(s):
// ramiframload_51 = (ramiframload_5 & (((always03 & LessThan1)) # (!\nRST~input_o )))

	.dataa(nRST),
	.datab(always03),
	.datac(LessThan1),
	.datad(ramiframload_5),
	.cin(gnd),
	.combout(ramiframload_51),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~9 .lut_mask = 16'hD500;
defparam \ramif.ramload[5]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N18
cycloneive_lcell_comb \ramif.ramload[6]~10 (
// Equation(s):
// ramiframload_6 = ((address_reg_a_0 & (ram_block3a381)) # (!address_reg_a_0 & ((ram_block3a64)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_6),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[6]~10 .lut_mask = 16'hD8FF;
defparam \ramif.ramload[6]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N28
cycloneive_lcell_comb \ramif.ramload[7]~11 (
// Equation(s):
// ramiframload_7 = ((address_reg_a_0 & (ram_block3a391)) # (!address_reg_a_0 & ((ram_block3a71)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_7),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[7]~11 .lut_mask = 16'hD8FF;
defparam \ramif.ramload[7]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N30
cycloneive_lcell_comb \ramif.ramload[8]~12 (
// Equation(s):
// ramiframload_8 = (always1 & ((address_reg_a_0 & (ram_block3a401)) # (!address_reg_a_0 & ((ram_block3a81)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_8),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[8]~12 .lut_mask = 16'h88C0;
defparam \ramif.ramload[8]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N8
cycloneive_lcell_comb \ramif.ramload[9]~13 (
// Equation(s):
// ramiframload_9 = ((address_reg_a_0 & ((ram_block3a412))) # (!address_reg_a_0 & (ram_block3a91))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_9),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[9]~13 .lut_mask = 16'hE4FF;
defparam \ramif.ramload[9]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N16
cycloneive_lcell_comb \ramif.ramload[10]~14 (
// Equation(s):
// ramiframload_10 = (always1 & ((address_reg_a_0 & (ram_block3a421)) # (!address_reg_a_0 & ((ram_block3a101)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_10),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[10]~14 .lut_mask = 16'hD800;
defparam \ramif.ramload[10]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N14
cycloneive_lcell_comb \ramif.ramload[11]~15 (
// Equation(s):
// ramiframload_11 = ((address_reg_a_0 & (ram_block3a431)) # (!address_reg_a_0 & ((ram_block3a112)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.cin(gnd),
	.combout(ramiframload_11),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[11]~15 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[11]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N18
cycloneive_lcell_comb \ramif.ramload[12]~16 (
// Equation(s):
// ramiframload_12 = ((address_reg_a_0 & ((ram_block3a441))) # (!address_reg_a_0 & (ram_block3a121))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.cin(gnd),
	.combout(ramiframload_12),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[12]~16 .lut_mask = 16'hFB73;
defparam \ramif.ramload[12]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N24
cycloneive_lcell_comb \ramif.ramload[13]~17 (
// Equation(s):
// ramiframload_13 = ((address_reg_a_0 & (ram_block3a451)) # (!address_reg_a_0 & ((ram_block3a131)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.cin(gnd),
	.combout(ramiframload_13),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[13]~17 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[13]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N12
cycloneive_lcell_comb \ramif.ramload[14]~18 (
// Equation(s):
// ramiframload_14 = (always1 & ((address_reg_a_0 & ((ram_block3a461))) # (!address_reg_a_0 & (ram_block3a141))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_14),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[14]~18 .lut_mask = 16'hE400;
defparam \ramif.ramload[14]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N6
cycloneive_lcell_comb \ramif.ramload[15]~19 (
// Equation(s):
// ramiframload_15 = ((address_reg_a_0 & (ram_block3a471)) # (!address_reg_a_0 & ((ram_block3a151)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.cin(gnd),
	.combout(ramiframload_15),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[15]~19 .lut_mask = 16'hBFB3;
defparam \ramif.ramload[15]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N0
cycloneive_lcell_comb \ramif.ramload[16]~20 (
// Equation(s):
// ramiframload_16 = (address_reg_a_0 & (ram_block3a481)) # (!address_reg_a_0 & ((ram_block3a161)))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.cin(gnd),
	.combout(ramiframload_16),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~20 .lut_mask = 16'hF3C0;
defparam \ramif.ramload[16]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N4
cycloneive_lcell_comb \ramif.ramload[16]~21 (
// Equation(s):
// ramiframload_161 = (ramiframload_16) # ((\nRST~input_o  & ((!LessThan1) # (!always03))))

	.dataa(nRST),
	.datab(always03),
	.datac(LessThan1),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(ramiframload_161),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~21 .lut_mask = 16'hFF2A;
defparam \ramif.ramload[16]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N6
cycloneive_lcell_comb \ramif.ramload[17]~22 (
// Equation(s):
// ramiframload_17 = (address_reg_a_0 & (ram_block3a491)) # (!address_reg_a_0 & ((ram_block3a171)))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.datad(gnd),
	.cin(gnd),
	.combout(ramiframload_17),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~22 .lut_mask = 16'hB8B8;
defparam \ramif.ramload[17]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N6
cycloneive_lcell_comb \ramif.ramload[17]~23 (
// Equation(s):
// ramiframload_171 = (ramiframload_17 & (((LessThan1 & always03)) # (!\nRST~input_o )))

	.dataa(ramiframload_17),
	.datab(nRST),
	.datac(LessThan1),
	.datad(always03),
	.cin(gnd),
	.combout(ramiframload_171),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~23 .lut_mask = 16'hA222;
defparam \ramif.ramload[17]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N28
cycloneive_lcell_comb \ramif.ramload[18]~24 (
// Equation(s):
// ramiframload_18 = (always1 & ((address_reg_a_0 & ((ram_block3a501))) # (!address_reg_a_0 & (ram_block3a181))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_18),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[18]~24 .lut_mask = 16'hE400;
defparam \ramif.ramload[18]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N24
cycloneive_lcell_comb \ramif.ramload[19]~25 (
// Equation(s):
// ramiframload_19 = (always1 & ((address_reg_a_0 & (ram_block3a512)) # (!address_reg_a_0 & ((ram_block3a191)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_19),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[19]~25 .lut_mask = 16'hA0C0;
defparam \ramif.ramload[19]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N14
cycloneive_lcell_comb \ramif.ramload[20]~26 (
// Equation(s):
// ramiframload_20 = ((address_reg_a_0 & (ram_block3a521)) # (!address_reg_a_0 & ((ram_block3a201)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.cin(gnd),
	.combout(ramiframload_20),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[20]~26 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[20]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N6
cycloneive_lcell_comb \ramif.ramload[21]~27 (
// Equation(s):
// ramiframload_211 = (always1 & ((address_reg_a_0 & ((ram_block3a531))) # (!address_reg_a_0 & (ram_block3a212))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_211),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[21]~27 .lut_mask = 16'hCA00;
defparam \ramif.ramload[21]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N0
cycloneive_lcell_comb \ramif.ramload[22]~28 (
// Equation(s):
// ramiframload_22 = ((address_reg_a_0 & (ram_block3a541)) # (!address_reg_a_0 & ((ram_block3a221)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_22),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[22]~28 .lut_mask = 16'hDDF5;
defparam \ramif.ramload[22]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N2
cycloneive_lcell_comb \ramif.ramload[23]~29 (
// Equation(s):
// ramiframload_23 = ((address_reg_a_0 & (ram_block3a551)) # (!address_reg_a_0 & ((ram_block3a231)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_23),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[23]~29 .lut_mask = 16'hB8FF;
defparam \ramif.ramload[23]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N20
cycloneive_lcell_comb \ramif.ramload[24]~30 (
// Equation(s):
// ramiframload_24 = (always1 & ((address_reg_a_0 & (ram_block3a561)) # (!address_reg_a_0 & ((ram_block3a241)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_24),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[24]~30 .lut_mask = 16'hD800;
defparam \ramif.ramload[24]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N0
cycloneive_lcell_comb \ramif.ramload[25]~31 (
// Equation(s):
// ramiframload_25 = ((address_reg_a_0 & ((ram_block3a571))) # (!address_reg_a_0 & (ram_block3a251))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.cin(gnd),
	.combout(ramiframload_25),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[25]~31 .lut_mask = 16'hFB73;
defparam \ramif.ramload[25]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N0
cycloneive_lcell_comb \ramif.ramload[26]~32 (
// Equation(s):
// ramiframload_26 = (address_reg_a_0 & ((ram_block3a581))) # (!address_reg_a_0 & (ram_block3a261))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.cin(gnd),
	.combout(ramiframload_26),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~32 .lut_mask = 16'hFC30;
defparam \ramif.ramload[26]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N18
cycloneive_lcell_comb \ramif.ramload[26]~33 (
// Equation(s):
// ramiframload_261 = (ramiframload_26 & (((always03 & LessThan1)) # (!\nRST~input_o )))

	.dataa(nRST),
	.datab(always03),
	.datac(LessThan1),
	.datad(ramiframload_26),
	.cin(gnd),
	.combout(ramiframload_261),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~33 .lut_mask = 16'hD500;
defparam \ramif.ramload[26]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N6
cycloneive_lcell_comb \ramif.ramload[27]~34 (
// Equation(s):
// ramiframload_27 = (address_reg_a_0 & (ram_block3a591)) # (!address_reg_a_0 & ((ram_block3a271)))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.cin(gnd),
	.combout(ramiframload_27),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~34 .lut_mask = 16'hF3C0;
defparam \ramif.ramload[27]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N24
cycloneive_lcell_comb \ramif.ramload[27]~35 (
// Equation(s):
// ramiframload_271 = (ramiframload_27) # ((\nRST~input_o  & ((!LessThan1) # (!always03))))

	.dataa(ramiframload_27),
	.datab(always03),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(ramiframload_271),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~35 .lut_mask = 16'hBFAA;
defparam \ramif.ramload[27]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N14
cycloneive_lcell_comb \ramif.ramload[28]~36 (
// Equation(s):
// ramiframload_28 = (address_reg_a_0 & (ram_block3a601)) # (!address_reg_a_0 & ((ram_block3a281)))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.cin(gnd),
	.combout(ramiframload_28),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~36 .lut_mask = 16'hF3C0;
defparam \ramif.ramload[28]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N6
cycloneive_lcell_comb \ramif.ramload[28]~37 (
// Equation(s):
// ramiframload_281 = (ramiframload_28) # ((\nRST~input_o  & ((!LessThan1) # (!always03))))

	.dataa(ramiframload_28),
	.datab(always03),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(ramiframload_281),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~37 .lut_mask = 16'hBFAA;
defparam \ramif.ramload[28]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N20
cycloneive_lcell_comb \ramif.ramload[29]~38 (
// Equation(s):
// ramiframload_29 = (address_reg_a_0 & (ram_block3a611)) # (!address_reg_a_0 & ((ram_block3a291)))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.datac(gnd),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.cin(gnd),
	.combout(ramiframload_29),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~38 .lut_mask = 16'hDD88;
defparam \ramif.ramload[29]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N8
cycloneive_lcell_comb \ramif.ramload[29]~39 (
// Equation(s):
// ramiframload_291 = (ramiframload_29) # ((\nRST~input_o  & ((!always03) # (!LessThan1))))

	.dataa(LessThan1),
	.datab(always03),
	.datac(nRST),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(ramiframload_291),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~39 .lut_mask = 16'hFF70;
defparam \ramif.ramload[29]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N30
cycloneive_lcell_comb \ramif.ramload[30]~40 (
// Equation(s):
// ramiframload_30 = (address_reg_a_0 & ((ram_block3a621))) # (!address_reg_a_0 & (ram_block3a301))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.cin(gnd),
	.combout(ramiframload_30),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~40 .lut_mask = 16'hFC30;
defparam \ramif.ramload[30]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N16
cycloneive_lcell_comb \ramif.ramload[30]~41 (
// Equation(s):
// ramiframload_301 = (ramiframload_30 & (((always03 & LessThan1)) # (!\nRST~input_o )))

	.dataa(nRST),
	.datab(always03),
	.datac(LessThan1),
	.datad(ramiframload_30),
	.cin(gnd),
	.combout(ramiframload_301),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~41 .lut_mask = 16'hD500;
defparam \ramif.ramload[30]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N12
cycloneive_lcell_comb \ramif.ramload[31]~42 (
// Equation(s):
// ramiframload_31 = (address_reg_a_0 & ((ram_block3a631))) # (!address_reg_a_0 & (ram_block3a312))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.cin(gnd),
	.combout(ramiframload_31),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~42 .lut_mask = 16'hFC30;
defparam \ramif.ramload[31]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N16
cycloneive_lcell_comb \ramif.ramload[31]~43 (
// Equation(s):
// ramiframload_311 = (ramiframload_31) # ((\nRST~input_o  & ((!LessThan1) # (!always03))))

	.dataa(always03),
	.datab(ramiframload_31),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(ramiframload_311),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~43 .lut_mask = 16'hDFCC;
defparam \ramif.ramload[31]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N7
dffeas \en[1] (
	.clk(CLK),
	.d(\ramif.ramREN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[1]),
	.prn(vcc));
// synopsys translate_off
defparam \en[1] .is_wysiwyg = "true";
defparam \en[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N29
dffeas \en[0] (
	.clk(CLK),
	.d(\ramif.ramWEN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[0]),
	.prn(vcc));
// synopsys translate_off
defparam \en[0] .is_wysiwyg = "true";
defparam \en[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N8
cycloneive_lcell_comb \always0~22 (
// Equation(s):
// \always0~22_combout  = (\ramREN~1_combout  & ((en[0] $ (\ramWEN~0_combout )) # (!en[1]))) # (!\ramREN~1_combout  & ((en[1]) # (en[0] $ (\ramWEN~0_combout ))))

	.dataa(\ramif.ramREN ),
	.datab(en[1]),
	.datac(en[0]),
	.datad(\ramif.ramWEN ),
	.cin(gnd),
	.combout(\always0~22_combout ),
	.cout());
// synopsys translate_off
defparam \always0~22 .lut_mask = 16'h6FF6;
defparam \always0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N22
cycloneive_lcell_comb \always0~23 (
// Equation(s):
// \always0~23_combout  = (((\always0~22_combout ) # (!always0)) # (!always01)) # (!always02)

	.dataa(always02),
	.datab(always01),
	.datac(\always0~22_combout ),
	.datad(always0),
	.cin(gnd),
	.combout(\always0~23_combout ),
	.cout());
// synopsys translate_off
defparam \always0~23 .lut_mask = 16'hF7FF;
defparam \always0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N12
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = (!\always0~23_combout  & (count[1] $ (((count[0] & !LessThan1)))))

	.dataa(count[0]),
	.datab(LessThan1),
	.datac(count[1]),
	.datad(\always0~23_combout ),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h00D2;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N13
dffeas \count[1] (
	.clk(CLK),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N22
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_combout  = (!count[1]) # (!count[0])

	.dataa(count[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(count[1]),
	.cin(gnd),
	.combout(\LessThan1~1_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h55FF;
defparam \LessThan1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N18
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = (!\always0~23_combout  & (count[2] $ (((!LessThan1 & !\LessThan1~1_combout )))))

	.dataa(\always0~23_combout ),
	.datab(LessThan1),
	.datac(count[2]),
	.datad(\LessThan1~1_combout ),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h5041;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N19
dffeas \count[2] (
	.clk(CLK),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N26
cycloneive_lcell_comb \count[0]~3 (
// Equation(s):
// \count[0]~3_combout  = (!\always0~23_combout  & (LessThan1 $ (!count[0])))

	.dataa(\always0~23_combout ),
	.datab(LessThan1),
	.datac(count[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \count[0]~3 .lut_mask = 16'h4141;
defparam \count[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N27
dffeas \count[0] (
	.clk(CLK),
	.d(\count[0]~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N28
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = (!\always0~23_combout  & count[3])

	.dataa(\always0~23_combout ),
	.datab(gnd),
	.datac(count[3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h5050;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N29
dffeas \count[3] (
	.clk(CLK),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N1
dffeas \addr[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr3),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[2] .is_wysiwyg = "true";
defparam \addr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N27
dffeas \addr[3] (
	.clk(CLK),
	.d(ramaddr2),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[3] .is_wysiwyg = "true";
defparam \addr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N0
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (\ramaddr~5_combout  & (addr[3] & (\ramaddr~7_combout  $ (!addr[2])))) # (!\ramaddr~5_combout  & (!addr[3] & (\ramaddr~7_combout  $ (!addr[2]))))

	.dataa(ramaddr2),
	.datab(ramaddr3),
	.datac(addr[2]),
	.datad(addr[3]),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'h8241;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N11
dffeas \addr[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[1] .is_wysiwyg = "true";
defparam \addr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N29
dffeas \addr[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[0] .is_wysiwyg = "true";
defparam \addr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N28
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (addr[1] & (\ramaddr~1_combout  & (addr[0] $ (!\ramaddr~3_combout )))) # (!addr[1] & (!\ramaddr~1_combout  & (addr[0] $ (!\ramaddr~3_combout ))))

	.dataa(addr[1]),
	.datab(ramaddr),
	.datac(addr[0]),
	.datad(ramaddr1),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h9009;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N14
cycloneive_lcell_comb \addr[5]~feeder (
// Equation(s):
// \addr[5]~feeder_combout  = \ramaddr~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(ramaddr4),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[5]~feeder .lut_mask = 16'hF0F0;
defparam \addr[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N15
dffeas \addr[5] (
	.clk(CLK),
	.d(\addr[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[5] .is_wysiwyg = "true";
defparam \addr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N1
dffeas \addr[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr5),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[4] .is_wysiwyg = "true";
defparam \addr[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N0
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// \always0~2_combout  = (\ramaddr~9_combout  & (addr[5] & (addr[4] $ (!\ramaddr~11_combout )))) # (!\ramaddr~9_combout  & (!addr[5] & (addr[4] $ (!\ramaddr~11_combout ))))

	.dataa(ramaddr4),
	.datab(addr[5]),
	.datac(addr[4]),
	.datad(ramaddr5),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'h9009;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N26
cycloneive_lcell_comb \addr[7]~feeder (
// Equation(s):
// \addr[7]~feeder_combout  = \ramaddr~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\addr[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[7]~feeder .lut_mask = 16'hFF00;
defparam \addr[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N27
dffeas \addr[7] (
	.clk(CLK),
	.d(\addr[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[7] .is_wysiwyg = "true";
defparam \addr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N9
dffeas \addr[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr7),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[6] .is_wysiwyg = "true";
defparam \addr[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N8
cycloneive_lcell_comb \always0~3 (
// Equation(s):
// \always0~3_combout  = (addr[7] & (\ramaddr~13_combout  & (\ramaddr~15_combout  $ (!addr[6])))) # (!addr[7] & (!\ramaddr~13_combout  & (\ramaddr~15_combout  $ (!addr[6]))))

	.dataa(addr[7]),
	.datab(ramaddr7),
	.datac(addr[6]),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\always0~3_combout ),
	.cout());
// synopsys translate_off
defparam \always0~3 .lut_mask = 16'h8241;
defparam \always0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N1
dffeas \addr[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr8),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[9] .is_wysiwyg = "true";
defparam \addr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N23
dffeas \addr[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr9),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[8] .is_wysiwyg = "true";
defparam \addr[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N22
cycloneive_lcell_comb \always0~5 (
// Equation(s):
// \always0~5_combout  = (addr[9] & (\ramaddr~17_combout  & (\ramaddr~19_combout  $ (!addr[8])))) # (!addr[9] & (!\ramaddr~17_combout  & (\ramaddr~19_combout  $ (!addr[8]))))

	.dataa(addr[9]),
	.datab(ramaddr9),
	.datac(addr[8]),
	.datad(ramaddr8),
	.cin(gnd),
	.combout(\always0~5_combout ),
	.cout());
// synopsys translate_off
defparam \always0~5 .lut_mask = 16'h8241;
defparam \always0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N27
dffeas \addr[15] (
	.clk(CLK),
	.d(ramaddr30),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[15] .is_wysiwyg = "true";
defparam \addr[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N21
dffeas \addr[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr15),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[14] .is_wysiwyg = "true";
defparam \addr[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N20
cycloneive_lcell_comb \always0~8 (
// Equation(s):
// \always0~8_combout  = (addr[15] & (!\ramaddr~29_combout  & (addr[14] $ (!\ramaddr~31_combout )))) # (!addr[15] & (\ramaddr~29_combout  & (addr[14] $ (!\ramaddr~31_combout ))))

	.dataa(addr[15]),
	.datab(ramaddr14),
	.datac(addr[14]),
	.datad(ramaddr15),
	.cin(gnd),
	.combout(\always0~8_combout ),
	.cout());
// synopsys translate_off
defparam \always0~8 .lut_mask = 16'h6006;
defparam \always0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N30
cycloneive_lcell_comb \addr[11]~feeder (
// Equation(s):
// \addr[11]~feeder_combout  = \ramaddr~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr10),
	.cin(gnd),
	.combout(\addr[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[11]~feeder .lut_mask = 16'hFF00;
defparam \addr[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N31
dffeas \addr[11] (
	.clk(CLK),
	.d(\addr[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[11] .is_wysiwyg = "true";
defparam \addr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N5
dffeas \addr[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr11),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[10] .is_wysiwyg = "true";
defparam \addr[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N4
cycloneive_lcell_comb \always0~6 (
// Equation(s):
// \always0~6_combout  = (\ramaddr~21_combout  & (addr[11] & (addr[10] $ (!\ramaddr~23_combout )))) # (!\ramaddr~21_combout  & (!addr[11] & (addr[10] $ (!\ramaddr~23_combout ))))

	.dataa(ramaddr10),
	.datab(addr[11]),
	.datac(addr[10]),
	.datad(ramaddr11),
	.cin(gnd),
	.combout(\always0~6_combout ),
	.cout());
// synopsys translate_off
defparam \always0~6 .lut_mask = 16'h9009;
defparam \always0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N6
cycloneive_lcell_comb \addr[13]~feeder (
// Equation(s):
// \addr[13]~feeder_combout  = \ramaddr~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr12),
	.cin(gnd),
	.combout(\addr[13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[13]~feeder .lut_mask = 16'hFF00;
defparam \addr[13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N7
dffeas \addr[13] (
	.clk(CLK),
	.d(\addr[13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[13] .is_wysiwyg = "true";
defparam \addr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N5
dffeas \addr[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr13),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[12] .is_wysiwyg = "true";
defparam \addr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N4
cycloneive_lcell_comb \always0~7 (
// Equation(s):
// \always0~7_combout  = (addr[13] & (\ramaddr~25_combout  & (\ramaddr~27_combout  $ (!addr[12])))) # (!addr[13] & (!\ramaddr~25_combout  & (\ramaddr~27_combout  $ (!addr[12]))))

	.dataa(addr[13]),
	.datab(ramaddr13),
	.datac(addr[12]),
	.datad(ramaddr12),
	.cin(gnd),
	.combout(\always0~7_combout ),
	.cout());
// synopsys translate_off
defparam \always0~7 .lut_mask = 16'h8241;
defparam \always0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N15
dffeas \addr[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr26),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[26] .is_wysiwyg = "true";
defparam \addr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N14
cycloneive_lcell_comb \always0~16 (
// Equation(s):
// \always0~16_combout  = (addr[27] & (\ramaddr~53_combout  & (\ramaddr~55_combout  $ (!addr[26])))) # (!addr[27] & (!\ramaddr~53_combout  & (\ramaddr~55_combout  $ (!addr[26]))))

	.dataa(addr[27]),
	.datab(ramaddr26),
	.datac(addr[26]),
	.datad(ramaddr25),
	.cin(gnd),
	.combout(\always0~16_combout ),
	.cout());
// synopsys translate_off
defparam \always0~16 .lut_mask = 16'h8241;
defparam \always0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N13
dffeas \addr[31] (
	.clk(CLK),
	.d(\ramif.ramaddr [31]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[31] .is_wysiwyg = "true";
defparam \addr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N23
dffeas \addr[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr29),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[30] .is_wysiwyg = "true";
defparam \addr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N22
cycloneive_lcell_comb \always0~18 (
// Equation(s):
// \always0~18_combout  = (\ramaddr~63_combout  & (addr[30] & (addr[31] $ (!\ramaddr~61_combout )))) # (!\ramaddr~63_combout  & (!addr[30] & (addr[31] $ (!\ramaddr~61_combout ))))

	.dataa(ramaddr29),
	.datab(addr[31]),
	.datac(addr[30]),
	.datad(\ramif.ramaddr [31]),
	.cin(gnd),
	.combout(\always0~18_combout ),
	.cout());
// synopsys translate_off
defparam \always0~18 .lut_mask = 16'h8421;
defparam \always0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N6
cycloneive_lcell_comb \addr[25]~feeder (
// Equation(s):
// \addr[25]~feeder_combout  = \ramaddr~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr23),
	.cin(gnd),
	.combout(\addr[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[25]~feeder .lut_mask = 16'hFF00;
defparam \addr[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N7
dffeas \addr[25] (
	.clk(CLK),
	.d(\addr[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[25] .is_wysiwyg = "true";
defparam \addr[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N29
dffeas \addr[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr24),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[24] .is_wysiwyg = "true";
defparam \addr[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N28
cycloneive_lcell_comb \always0~15 (
// Equation(s):
// \always0~15_combout  = (\ramaddr~51_combout  & (addr[24] & (addr[25] $ (!\ramaddr~49_combout )))) # (!\ramaddr~51_combout  & (!addr[24] & (addr[25] $ (!\ramaddr~49_combout ))))

	.dataa(ramaddr24),
	.datab(addr[25]),
	.datac(addr[24]),
	.datad(ramaddr23),
	.cin(gnd),
	.combout(\always0~15_combout ),
	.cout());
// synopsys translate_off
defparam \always0~15 .lut_mask = 16'h8421;
defparam \always0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N5
dffeas \addr[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr28),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[28] .is_wysiwyg = "true";
defparam \addr[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N4
cycloneive_lcell_comb \always0~17 (
// Equation(s):
// \always0~17_combout  = (addr[29] & (\ramaddr~57_combout  & (addr[28] $ (!\ramaddr~59_combout )))) # (!addr[29] & (!\ramaddr~57_combout  & (addr[28] $ (!\ramaddr~59_combout ))))

	.dataa(addr[29]),
	.datab(ramaddr27),
	.datac(addr[28]),
	.datad(ramaddr28),
	.cin(gnd),
	.combout(\always0~17_combout ),
	.cout());
// synopsys translate_off
defparam \always0~17 .lut_mask = 16'h9009;
defparam \always0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N8
cycloneive_lcell_comb \always0~19 (
// Equation(s):
// \always0~19_combout  = (\always0~16_combout  & (\always0~18_combout  & (\always0~15_combout  & \always0~17_combout )))

	.dataa(\always0~16_combout ),
	.datab(\always0~18_combout ),
	.datac(\always0~15_combout ),
	.datad(\always0~17_combout ),
	.cin(gnd),
	.combout(\always0~19_combout ),
	.cout());
// synopsys translate_off
defparam \always0~19 .lut_mask = 16'h8000;
defparam \always0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N7
dffeas \addr[19] (
	.clk(CLK),
	.d(\ramif.ramaddr [19]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[19] .is_wysiwyg = "true";
defparam \addr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N21
dffeas \addr[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr18),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[18] .is_wysiwyg = "true";
defparam \addr[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N20
cycloneive_lcell_comb \always0~11 (
// Equation(s):
// \always0~11_combout  = (\ramaddr~37_combout  & (addr[19] & (addr[18] $ (!\ramaddr~39_combout )))) # (!\ramaddr~37_combout  & (!addr[19] & (addr[18] $ (!\ramaddr~39_combout ))))

	.dataa(\ramif.ramaddr [19]),
	.datab(addr[19]),
	.datac(addr[18]),
	.datad(ramaddr18),
	.cin(gnd),
	.combout(\always0~11_combout ),
	.cout());
// synopsys translate_off
defparam \always0~11 .lut_mask = 16'h9009;
defparam \always0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N17
dffeas \addr[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr20),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[20] .is_wysiwyg = "true";
defparam \addr[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N16
cycloneive_lcell_comb \always0~12 (
// Equation(s):
// \always0~12_combout  = (addr[21] & (\ramaddr~41_combout  & (\ramaddr~43_combout  $ (!addr[20])))) # (!addr[21] & (!\ramaddr~41_combout  & (\ramaddr~43_combout  $ (!addr[20]))))

	.dataa(addr[21]),
	.datab(ramaddr20),
	.datac(addr[20]),
	.datad(ramaddr19),
	.cin(gnd),
	.combout(\always0~12_combout ),
	.cout());
// synopsys translate_off
defparam \always0~12 .lut_mask = 16'h8241;
defparam \always0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N25
dffeas \addr[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr17),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[16] .is_wysiwyg = "true";
defparam \addr[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N24
cycloneive_lcell_comb \always0~10 (
// Equation(s):
// \always0~10_combout  = (addr[17] & (\ramaddr~33_combout  & (addr[16] $ (!\ramaddr~35_combout )))) # (!addr[17] & (!\ramaddr~33_combout  & (addr[16] $ (!\ramaddr~35_combout ))))

	.dataa(addr[17]),
	.datab(ramaddr16),
	.datac(addr[16]),
	.datad(ramaddr17),
	.cin(gnd),
	.combout(\always0~10_combout ),
	.cout());
// synopsys translate_off
defparam \always0~10 .lut_mask = 16'h9009;
defparam \always0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y43_N17
dffeas \addr[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr22),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[22] .is_wysiwyg = "true";
defparam \addr[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N16
cycloneive_lcell_comb \always0~13 (
// Equation(s):
// \always0~13_combout  = (addr[23] & (\ramaddr~45_combout  & (\ramaddr~47_combout  $ (!addr[22])))) # (!addr[23] & (!\ramaddr~45_combout  & (\ramaddr~47_combout  $ (!addr[22]))))

	.dataa(addr[23]),
	.datab(ramaddr22),
	.datac(addr[22]),
	.datad(ramaddr21),
	.cin(gnd),
	.combout(\always0~13_combout ),
	.cout());
// synopsys translate_off
defparam \always0~13 .lut_mask = 16'h8241;
defparam \always0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N10
cycloneive_lcell_comb \always0~14 (
// Equation(s):
// \always0~14_combout  = (\always0~11_combout  & (\always0~12_combout  & (\always0~10_combout  & \always0~13_combout )))

	.dataa(\always0~11_combout ),
	.datab(\always0~12_combout ),
	.datac(\always0~10_combout ),
	.datad(\always0~13_combout ),
	.cin(gnd),
	.combout(\always0~14_combout ),
	.cout());
// synopsys translate_off
defparam \always0~14 .lut_mask = 16'h8000;
defparam \always0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N12
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// \always1~0_combout  = (LessThan1 & always01)

	.dataa(gnd),
	.datab(gnd),
	.datac(LessThan1),
	.datad(always01),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'hF000;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module altsyncram_1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



altsyncram_99f1 auto_generated(
	.ram_block3a32(ram_block3a32),
	.ram_block3a0(ram_block3a0),
	.ram_block3a33(ram_block3a33),
	.ram_block3a1(ram_block3a1),
	.ram_block3a34(ram_block3a34),
	.ram_block3a2(ram_block3a2),
	.ram_block3a35(ram_block3a35),
	.ram_block3a3(ram_block3a3),
	.ram_block3a36(ram_block3a36),
	.ram_block3a4(ram_block3a4),
	.ram_block3a37(ram_block3a37),
	.ram_block3a5(ram_block3a5),
	.ram_block3a38(ram_block3a38),
	.ram_block3a6(ram_block3a6),
	.ram_block3a39(ram_block3a39),
	.ram_block3a7(ram_block3a7),
	.ram_block3a40(ram_block3a40),
	.ram_block3a8(ram_block3a8),
	.ram_block3a41(ram_block3a41),
	.ram_block3a9(ram_block3a9),
	.ram_block3a42(ram_block3a42),
	.ram_block3a10(ram_block3a10),
	.ram_block3a43(ram_block3a43),
	.ram_block3a11(ram_block3a11),
	.ram_block3a44(ram_block3a44),
	.ram_block3a12(ram_block3a12),
	.ram_block3a45(ram_block3a45),
	.ram_block3a13(ram_block3a13),
	.ram_block3a46(ram_block3a46),
	.ram_block3a14(ram_block3a14),
	.ram_block3a47(ram_block3a47),
	.ram_block3a15(ram_block3a15),
	.ram_block3a48(ram_block3a48),
	.ram_block3a16(ram_block3a16),
	.ram_block3a49(ram_block3a49),
	.ram_block3a17(ram_block3a17),
	.ram_block3a50(ram_block3a50),
	.ram_block3a18(ram_block3a18),
	.ram_block3a51(ram_block3a51),
	.ram_block3a19(ram_block3a19),
	.ram_block3a52(ram_block3a52),
	.ram_block3a20(ram_block3a20),
	.ram_block3a53(ram_block3a53),
	.ram_block3a21(ram_block3a21),
	.ram_block3a54(ram_block3a54),
	.ram_block3a22(ram_block3a22),
	.ram_block3a55(ram_block3a55),
	.ram_block3a23(ram_block3a23),
	.ram_block3a56(ram_block3a56),
	.ram_block3a24(ram_block3a24),
	.ram_block3a57(ram_block3a57),
	.ram_block3a25(ram_block3a25),
	.ram_block3a58(ram_block3a58),
	.ram_block3a26(ram_block3a26),
	.ram_block3a59(ram_block3a59),
	.ram_block3a27(ram_block3a27),
	.ram_block3a60(ram_block3a60),
	.ram_block3a28(ram_block3a28),
	.ram_block3a61(ram_block3a61),
	.ram_block3a29(ram_block3a29),
	.ram_block3a62(ram_block3a62),
	.ram_block3a30(ram_block3a30),
	.ram_block3a63(ram_block3a63),
	.ram_block3a31(ram_block3a31),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.ramaddr1(ramaddr1),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_99f1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram1|ram_block3a32~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a0~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a33~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a1~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a34~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a2~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a35~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a3~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a36~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a4~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a37~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a5~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a38~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a6~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a39~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a7~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a40~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a8~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a41~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a9~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a42~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a10~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a43~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a11~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a44~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a12~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a45~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a13~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a46~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a14~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a47~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a15~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a48~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a16~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a49~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a17~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a50~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a18~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a51~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a19~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a52~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a20~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a53~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a21~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a54~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a22~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a55~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a23~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a56~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a24~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a57~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a25~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a58~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a26~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a59~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a27~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a60~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a28~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a61~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a29~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a62~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a30~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a63~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a31~PORTBDATAOUT0 ;
wire \mgl_prim2|sdr~0_combout ;
wire [0:0] \altsyncram1|address_reg_b ;
wire [31:0] \mgl_prim2|ram_rom_data_reg ;
wire [13:0] \mgl_prim2|ram_rom_addr_reg ;


sld_mod_ram_rom mgl_prim2(
	.ram_block3a32(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a0(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a33(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a1(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a34(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a2(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a35(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a3(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a36(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a4(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a37(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a5(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a38(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a6(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a39(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a7(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a40(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a8(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a41(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a9(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a42(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a10(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a43(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a11(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a44(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a12(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a45(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a13(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a46(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a14(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a47(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a15(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a48(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a16(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a49(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a17(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a50(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a18(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a51(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a19(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a52(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a20(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a53(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a21(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a54(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a22(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a55(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a23(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a56(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a24(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a57(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a25(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a58(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a26(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a59(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a27(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a60(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a28(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a61(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a29(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a62(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a30(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a63(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a31(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.is_in_use_reg1(is_in_use_reg),
	.ram_rom_data_reg_0(\mgl_prim2|ram_rom_data_reg [0]),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.ram_rom_addr_reg_0(\mgl_prim2|ram_rom_addr_reg [0]),
	.ram_rom_addr_reg_1(\mgl_prim2|ram_rom_addr_reg [1]),
	.ram_rom_addr_reg_2(\mgl_prim2|ram_rom_addr_reg [2]),
	.ram_rom_addr_reg_3(\mgl_prim2|ram_rom_addr_reg [3]),
	.ram_rom_addr_reg_4(\mgl_prim2|ram_rom_addr_reg [4]),
	.ram_rom_addr_reg_5(\mgl_prim2|ram_rom_addr_reg [5]),
	.ram_rom_addr_reg_6(\mgl_prim2|ram_rom_addr_reg [6]),
	.ram_rom_addr_reg_7(\mgl_prim2|ram_rom_addr_reg [7]),
	.ram_rom_addr_reg_8(\mgl_prim2|ram_rom_addr_reg [8]),
	.ram_rom_addr_reg_9(\mgl_prim2|ram_rom_addr_reg [9]),
	.ram_rom_addr_reg_10(\mgl_prim2|ram_rom_addr_reg [10]),
	.ram_rom_addr_reg_11(\mgl_prim2|ram_rom_addr_reg [11]),
	.ram_rom_addr_reg_12(\mgl_prim2|ram_rom_addr_reg [12]),
	.ram_rom_data_reg_1(\mgl_prim2|ram_rom_data_reg [1]),
	.ram_rom_data_reg_2(\mgl_prim2|ram_rom_data_reg [2]),
	.ram_rom_data_reg_3(\mgl_prim2|ram_rom_data_reg [3]),
	.ram_rom_data_reg_4(\mgl_prim2|ram_rom_data_reg [4]),
	.ram_rom_data_reg_5(\mgl_prim2|ram_rom_data_reg [5]),
	.ram_rom_data_reg_6(\mgl_prim2|ram_rom_data_reg [6]),
	.ram_rom_data_reg_7(\mgl_prim2|ram_rom_data_reg [7]),
	.ram_rom_data_reg_8(\mgl_prim2|ram_rom_data_reg [8]),
	.ram_rom_data_reg_9(\mgl_prim2|ram_rom_data_reg [9]),
	.ram_rom_data_reg_10(\mgl_prim2|ram_rom_data_reg [10]),
	.ram_rom_data_reg_11(\mgl_prim2|ram_rom_data_reg [11]),
	.ram_rom_data_reg_12(\mgl_prim2|ram_rom_data_reg [12]),
	.ram_rom_data_reg_13(\mgl_prim2|ram_rom_data_reg [13]),
	.ram_rom_data_reg_14(\mgl_prim2|ram_rom_data_reg [14]),
	.ram_rom_data_reg_15(\mgl_prim2|ram_rom_data_reg [15]),
	.ram_rom_data_reg_16(\mgl_prim2|ram_rom_data_reg [16]),
	.ram_rom_data_reg_17(\mgl_prim2|ram_rom_data_reg [17]),
	.ram_rom_data_reg_18(\mgl_prim2|ram_rom_data_reg [18]),
	.ram_rom_data_reg_19(\mgl_prim2|ram_rom_data_reg [19]),
	.ram_rom_data_reg_20(\mgl_prim2|ram_rom_data_reg [20]),
	.ram_rom_data_reg_21(\mgl_prim2|ram_rom_data_reg [21]),
	.ram_rom_data_reg_22(\mgl_prim2|ram_rom_data_reg [22]),
	.ram_rom_data_reg_23(\mgl_prim2|ram_rom_data_reg [23]),
	.ram_rom_data_reg_24(\mgl_prim2|ram_rom_data_reg [24]),
	.ram_rom_data_reg_25(\mgl_prim2|ram_rom_data_reg [25]),
	.ram_rom_data_reg_26(\mgl_prim2|ram_rom_data_reg [26]),
	.ram_rom_data_reg_27(\mgl_prim2|ram_rom_data_reg [27]),
	.ram_rom_data_reg_28(\mgl_prim2|ram_rom_data_reg [28]),
	.ram_rom_data_reg_29(\mgl_prim2|ram_rom_data_reg [29]),
	.ram_rom_data_reg_30(\mgl_prim2|ram_rom_data_reg [30]),
	.ram_rom_data_reg_31(\mgl_prim2|ram_rom_data_reg [31]),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.ir_in({gnd,irf_reg_3_1,gnd,gnd,irf_reg_0_1}),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.raw_tck(altera_internal_jtag1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

altsyncram_fta2 altsyncram1(
	.ram_block3a321(ram_block3a32),
	.ram_block3a322(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a01(ram_block3a0),
	.ram_block3a02(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a331(ram_block3a33),
	.ram_block3a332(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a110(ram_block3a1),
	.ram_block3a111(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a341(ram_block3a34),
	.ram_block3a342(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a210(ram_block3a2),
	.ram_block3a211(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a351(ram_block3a35),
	.ram_block3a352(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a310(ram_block3a3),
	.ram_block3a311(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a361(ram_block3a36),
	.ram_block3a362(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a410(ram_block3a4),
	.ram_block3a411(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a371(ram_block3a37),
	.ram_block3a372(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a510(ram_block3a5),
	.ram_block3a511(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a381(ram_block3a38),
	.ram_block3a382(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a64(ram_block3a6),
	.ram_block3a65(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a391(ram_block3a39),
	.ram_block3a392(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a71(ram_block3a7),
	.ram_block3a72(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a401(ram_block3a40),
	.ram_block3a402(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a81(ram_block3a8),
	.ram_block3a82(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a412(ram_block3a41),
	.ram_block3a413(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a91(ram_block3a9),
	.ram_block3a92(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a421(ram_block3a42),
	.ram_block3a422(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a101(ram_block3a10),
	.ram_block3a102(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a431(ram_block3a43),
	.ram_block3a432(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a112(ram_block3a11),
	.ram_block3a113(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a441(ram_block3a44),
	.ram_block3a442(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a121(ram_block3a12),
	.ram_block3a122(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a451(ram_block3a45),
	.ram_block3a452(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a131(ram_block3a13),
	.ram_block3a132(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a461(ram_block3a46),
	.ram_block3a462(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a141(ram_block3a14),
	.ram_block3a142(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a471(ram_block3a47),
	.ram_block3a472(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a151(ram_block3a15),
	.ram_block3a152(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a481(ram_block3a48),
	.ram_block3a482(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a161(ram_block3a16),
	.ram_block3a162(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a491(ram_block3a49),
	.ram_block3a492(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a171(ram_block3a17),
	.ram_block3a172(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a501(ram_block3a50),
	.ram_block3a502(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a181(ram_block3a18),
	.ram_block3a182(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a512(ram_block3a51),
	.ram_block3a513(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a191(ram_block3a19),
	.ram_block3a192(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a521(ram_block3a52),
	.ram_block3a522(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a201(ram_block3a20),
	.ram_block3a202(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a531(ram_block3a53),
	.ram_block3a532(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a212(ram_block3a21),
	.ram_block3a213(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a541(ram_block3a54),
	.ram_block3a542(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a221(ram_block3a22),
	.ram_block3a222(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a551(ram_block3a55),
	.ram_block3a552(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a231(ram_block3a23),
	.ram_block3a232(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a561(ram_block3a56),
	.ram_block3a562(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a241(ram_block3a24),
	.ram_block3a242(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a571(ram_block3a57),
	.ram_block3a572(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a251(ram_block3a25),
	.ram_block3a252(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a581(ram_block3a58),
	.ram_block3a582(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a261(ram_block3a26),
	.ram_block3a262(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a591(ram_block3a59),
	.ram_block3a592(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a271(ram_block3a27),
	.ram_block3a272(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a601(ram_block3a60),
	.ram_block3a602(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a281(ram_block3a28),
	.ram_block3a282(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a611(ram_block3a61),
	.ram_block3a612(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a291(ram_block3a29),
	.ram_block3a292(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a621(ram_block3a62),
	.ram_block3a622(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a301(ram_block3a30),
	.ram_block3a302(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a631(ram_block3a63),
	.ram_block3a632(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a312(ram_block3a31),
	.ram_block3a313(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.data_b({\mgl_prim2|ram_rom_data_reg [31],\mgl_prim2|ram_rom_data_reg [30],\mgl_prim2|ram_rom_data_reg [29],\mgl_prim2|ram_rom_data_reg [28],\mgl_prim2|ram_rom_data_reg [27],\mgl_prim2|ram_rom_data_reg [26],\mgl_prim2|ram_rom_data_reg [25],\mgl_prim2|ram_rom_data_reg [24],\mgl_prim2|ram_rom_data_reg [23],
\mgl_prim2|ram_rom_data_reg [22],\mgl_prim2|ram_rom_data_reg [21],\mgl_prim2|ram_rom_data_reg [20],\mgl_prim2|ram_rom_data_reg [19],\mgl_prim2|ram_rom_data_reg [18],\mgl_prim2|ram_rom_data_reg [17],\mgl_prim2|ram_rom_data_reg [16],\mgl_prim2|ram_rom_data_reg [15],\mgl_prim2|ram_rom_data_reg [14],
\mgl_prim2|ram_rom_data_reg [13],\mgl_prim2|ram_rom_data_reg [12],\mgl_prim2|ram_rom_data_reg [11],\mgl_prim2|ram_rom_data_reg [10],\mgl_prim2|ram_rom_data_reg [9],\mgl_prim2|ram_rom_data_reg [8],\mgl_prim2|ram_rom_data_reg [7],\mgl_prim2|ram_rom_data_reg [6],\mgl_prim2|ram_rom_data_reg [5],
\mgl_prim2|ram_rom_data_reg [4],\mgl_prim2|ram_rom_data_reg [3],\mgl_prim2|ram_rom_data_reg [2],\mgl_prim2|ram_rom_data_reg [1],\mgl_prim2|ram_rom_data_reg [0]}),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.address_b({gnd,\mgl_prim2|ram_rom_addr_reg [12],\mgl_prim2|ram_rom_addr_reg [11],\mgl_prim2|ram_rom_addr_reg [10],\mgl_prim2|ram_rom_addr_reg [9],\mgl_prim2|ram_rom_addr_reg [8],\mgl_prim2|ram_rom_addr_reg [7],\mgl_prim2|ram_rom_addr_reg [6],\mgl_prim2|ram_rom_addr_reg [5],\mgl_prim2|ram_rom_addr_reg [4],
\mgl_prim2|ram_rom_addr_reg [3],\mgl_prim2|ram_rom_addr_reg [2],\mgl_prim2|ram_rom_addr_reg [1],\mgl_prim2|ram_rom_addr_reg [0]}),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.ramaddr1(ramaddr1),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.clock1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_fta2 (
	ram_block3a321,
	ram_block3a322,
	ram_block3a01,
	ram_block3a02,
	ram_block3a331,
	ram_block3a332,
	ram_block3a110,
	ram_block3a111,
	ram_block3a341,
	ram_block3a342,
	ram_block3a210,
	ram_block3a211,
	ram_block3a351,
	ram_block3a352,
	ram_block3a310,
	ram_block3a311,
	ram_block3a361,
	ram_block3a362,
	ram_block3a410,
	ram_block3a411,
	ram_block3a371,
	ram_block3a372,
	ram_block3a510,
	ram_block3a511,
	ram_block3a381,
	ram_block3a382,
	ram_block3a64,
	ram_block3a65,
	ram_block3a391,
	ram_block3a392,
	ram_block3a71,
	ram_block3a72,
	ram_block3a401,
	ram_block3a402,
	ram_block3a81,
	ram_block3a82,
	ram_block3a412,
	ram_block3a413,
	ram_block3a91,
	ram_block3a92,
	ram_block3a421,
	ram_block3a422,
	ram_block3a101,
	ram_block3a102,
	ram_block3a431,
	ram_block3a432,
	ram_block3a112,
	ram_block3a113,
	ram_block3a441,
	ram_block3a442,
	ram_block3a121,
	ram_block3a122,
	ram_block3a451,
	ram_block3a452,
	ram_block3a131,
	ram_block3a132,
	ram_block3a461,
	ram_block3a462,
	ram_block3a141,
	ram_block3a142,
	ram_block3a471,
	ram_block3a472,
	ram_block3a151,
	ram_block3a152,
	ram_block3a481,
	ram_block3a482,
	ram_block3a161,
	ram_block3a162,
	ram_block3a491,
	ram_block3a492,
	ram_block3a171,
	ram_block3a172,
	ram_block3a501,
	ram_block3a502,
	ram_block3a181,
	ram_block3a182,
	ram_block3a512,
	ram_block3a513,
	ram_block3a191,
	ram_block3a192,
	ram_block3a521,
	ram_block3a522,
	ram_block3a201,
	ram_block3a202,
	ram_block3a531,
	ram_block3a532,
	ram_block3a212,
	ram_block3a213,
	ram_block3a541,
	ram_block3a542,
	ram_block3a221,
	ram_block3a222,
	ram_block3a551,
	ram_block3a552,
	ram_block3a231,
	ram_block3a232,
	ram_block3a561,
	ram_block3a562,
	ram_block3a241,
	ram_block3a242,
	ram_block3a571,
	ram_block3a572,
	ram_block3a251,
	ram_block3a252,
	ram_block3a581,
	ram_block3a582,
	ram_block3a261,
	ram_block3a262,
	ram_block3a591,
	ram_block3a592,
	ram_block3a271,
	ram_block3a272,
	ram_block3a601,
	ram_block3a602,
	ram_block3a281,
	ram_block3a282,
	ram_block3a611,
	ram_block3a612,
	ram_block3a291,
	ram_block3a292,
	ram_block3a621,
	ram_block3a622,
	ram_block3a301,
	ram_block3a302,
	ram_block3a631,
	ram_block3a632,
	ram_block3a312,
	ram_block3a313,
	data_b,
	ram_rom_addr_reg_13,
	address_b,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	sdr,
	data_a,
	address_reg_b_0,
	ramaddr1,
	irf_reg_2_1,
	state_5,
	clock1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a321;
output 	ram_block3a322;
output 	ram_block3a01;
output 	ram_block3a02;
output 	ram_block3a331;
output 	ram_block3a332;
output 	ram_block3a110;
output 	ram_block3a111;
output 	ram_block3a341;
output 	ram_block3a342;
output 	ram_block3a210;
output 	ram_block3a211;
output 	ram_block3a351;
output 	ram_block3a352;
output 	ram_block3a310;
output 	ram_block3a311;
output 	ram_block3a361;
output 	ram_block3a362;
output 	ram_block3a410;
output 	ram_block3a411;
output 	ram_block3a371;
output 	ram_block3a372;
output 	ram_block3a510;
output 	ram_block3a511;
output 	ram_block3a381;
output 	ram_block3a382;
output 	ram_block3a64;
output 	ram_block3a65;
output 	ram_block3a391;
output 	ram_block3a392;
output 	ram_block3a71;
output 	ram_block3a72;
output 	ram_block3a401;
output 	ram_block3a402;
output 	ram_block3a81;
output 	ram_block3a82;
output 	ram_block3a412;
output 	ram_block3a413;
output 	ram_block3a91;
output 	ram_block3a92;
output 	ram_block3a421;
output 	ram_block3a422;
output 	ram_block3a101;
output 	ram_block3a102;
output 	ram_block3a431;
output 	ram_block3a432;
output 	ram_block3a112;
output 	ram_block3a113;
output 	ram_block3a441;
output 	ram_block3a442;
output 	ram_block3a121;
output 	ram_block3a122;
output 	ram_block3a451;
output 	ram_block3a452;
output 	ram_block3a131;
output 	ram_block3a132;
output 	ram_block3a461;
output 	ram_block3a462;
output 	ram_block3a141;
output 	ram_block3a142;
output 	ram_block3a471;
output 	ram_block3a472;
output 	ram_block3a151;
output 	ram_block3a152;
output 	ram_block3a481;
output 	ram_block3a482;
output 	ram_block3a161;
output 	ram_block3a162;
output 	ram_block3a491;
output 	ram_block3a492;
output 	ram_block3a171;
output 	ram_block3a172;
output 	ram_block3a501;
output 	ram_block3a502;
output 	ram_block3a181;
output 	ram_block3a182;
output 	ram_block3a512;
output 	ram_block3a513;
output 	ram_block3a191;
output 	ram_block3a192;
output 	ram_block3a521;
output 	ram_block3a522;
output 	ram_block3a201;
output 	ram_block3a202;
output 	ram_block3a531;
output 	ram_block3a532;
output 	ram_block3a212;
output 	ram_block3a213;
output 	ram_block3a541;
output 	ram_block3a542;
output 	ram_block3a221;
output 	ram_block3a222;
output 	ram_block3a551;
output 	ram_block3a552;
output 	ram_block3a231;
output 	ram_block3a232;
output 	ram_block3a561;
output 	ram_block3a562;
output 	ram_block3a241;
output 	ram_block3a242;
output 	ram_block3a571;
output 	ram_block3a572;
output 	ram_block3a251;
output 	ram_block3a252;
output 	ram_block3a581;
output 	ram_block3a582;
output 	ram_block3a261;
output 	ram_block3a262;
output 	ram_block3a591;
output 	ram_block3a592;
output 	ram_block3a271;
output 	ram_block3a272;
output 	ram_block3a601;
output 	ram_block3a602;
output 	ram_block3a281;
output 	ram_block3a282;
output 	ram_block3a611;
output 	ram_block3a612;
output 	ram_block3a291;
output 	ram_block3a292;
output 	ram_block3a621;
output 	ram_block3a622;
output 	ram_block3a301;
output 	ram_block3a302;
output 	ram_block3a631;
output 	ram_block3a632;
output 	ram_block3a312;
output 	ram_block3a313;
input 	[31:0] data_b;
input 	ram_rom_addr_reg_13;
input 	[13:0] address_b;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
input 	sdr;
input 	[31:0] data_a;
output 	address_reg_b_0;
input 	ramaddr1;
input 	irf_reg_2_1;
input 	state_5;
input 	clock1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \decode4|eq_node[1]~0_combout ;
wire \decode5|eq_node[1]~0_combout ;
wire \decode4|eq_node[0]~1_combout ;
wire \decode5|eq_node[0]~1_combout ;
wire \address_reg_b[0]~feeder_combout ;

wire [0:0] ram_block3a32_PORTADATAOUT_bus;
wire [0:0] ram_block3a32_PORTBDATAOUT_bus;
wire [0:0] ram_block3a0_PORTADATAOUT_bus;
wire [0:0] ram_block3a0_PORTBDATAOUT_bus;
wire [0:0] ram_block3a33_PORTADATAOUT_bus;
wire [0:0] ram_block3a33_PORTBDATAOUT_bus;
wire [0:0] ram_block3a1_PORTADATAOUT_bus;
wire [0:0] ram_block3a1_PORTBDATAOUT_bus;
wire [0:0] ram_block3a34_PORTADATAOUT_bus;
wire [0:0] ram_block3a34_PORTBDATAOUT_bus;
wire [0:0] ram_block3a2_PORTADATAOUT_bus;
wire [0:0] ram_block3a2_PORTBDATAOUT_bus;
wire [0:0] ram_block3a35_PORTADATAOUT_bus;
wire [0:0] ram_block3a35_PORTBDATAOUT_bus;
wire [0:0] ram_block3a3_PORTADATAOUT_bus;
wire [0:0] ram_block3a3_PORTBDATAOUT_bus;
wire [0:0] ram_block3a36_PORTADATAOUT_bus;
wire [0:0] ram_block3a36_PORTBDATAOUT_bus;
wire [0:0] ram_block3a4_PORTADATAOUT_bus;
wire [0:0] ram_block3a4_PORTBDATAOUT_bus;
wire [0:0] ram_block3a37_PORTADATAOUT_bus;
wire [0:0] ram_block3a37_PORTBDATAOUT_bus;
wire [0:0] ram_block3a5_PORTADATAOUT_bus;
wire [0:0] ram_block3a5_PORTBDATAOUT_bus;
wire [0:0] ram_block3a38_PORTADATAOUT_bus;
wire [0:0] ram_block3a38_PORTBDATAOUT_bus;
wire [0:0] ram_block3a6_PORTADATAOUT_bus;
wire [0:0] ram_block3a6_PORTBDATAOUT_bus;
wire [0:0] ram_block3a39_PORTADATAOUT_bus;
wire [0:0] ram_block3a39_PORTBDATAOUT_bus;
wire [0:0] ram_block3a7_PORTADATAOUT_bus;
wire [0:0] ram_block3a7_PORTBDATAOUT_bus;
wire [0:0] ram_block3a40_PORTADATAOUT_bus;
wire [0:0] ram_block3a40_PORTBDATAOUT_bus;
wire [0:0] ram_block3a8_PORTADATAOUT_bus;
wire [0:0] ram_block3a8_PORTBDATAOUT_bus;
wire [0:0] ram_block3a41_PORTADATAOUT_bus;
wire [0:0] ram_block3a41_PORTBDATAOUT_bus;
wire [0:0] ram_block3a9_PORTADATAOUT_bus;
wire [0:0] ram_block3a9_PORTBDATAOUT_bus;
wire [0:0] ram_block3a42_PORTADATAOUT_bus;
wire [0:0] ram_block3a42_PORTBDATAOUT_bus;
wire [0:0] ram_block3a10_PORTADATAOUT_bus;
wire [0:0] ram_block3a10_PORTBDATAOUT_bus;
wire [0:0] ram_block3a43_PORTADATAOUT_bus;
wire [0:0] ram_block3a43_PORTBDATAOUT_bus;
wire [0:0] ram_block3a11_PORTADATAOUT_bus;
wire [0:0] ram_block3a11_PORTBDATAOUT_bus;
wire [0:0] ram_block3a44_PORTADATAOUT_bus;
wire [0:0] ram_block3a44_PORTBDATAOUT_bus;
wire [0:0] ram_block3a12_PORTADATAOUT_bus;
wire [0:0] ram_block3a12_PORTBDATAOUT_bus;
wire [0:0] ram_block3a45_PORTADATAOUT_bus;
wire [0:0] ram_block3a45_PORTBDATAOUT_bus;
wire [0:0] ram_block3a13_PORTADATAOUT_bus;
wire [0:0] ram_block3a13_PORTBDATAOUT_bus;
wire [0:0] ram_block3a46_PORTADATAOUT_bus;
wire [0:0] ram_block3a46_PORTBDATAOUT_bus;
wire [0:0] ram_block3a14_PORTADATAOUT_bus;
wire [0:0] ram_block3a14_PORTBDATAOUT_bus;
wire [0:0] ram_block3a47_PORTADATAOUT_bus;
wire [0:0] ram_block3a47_PORTBDATAOUT_bus;
wire [0:0] ram_block3a15_PORTADATAOUT_bus;
wire [0:0] ram_block3a15_PORTBDATAOUT_bus;
wire [0:0] ram_block3a48_PORTADATAOUT_bus;
wire [0:0] ram_block3a48_PORTBDATAOUT_bus;
wire [0:0] ram_block3a16_PORTADATAOUT_bus;
wire [0:0] ram_block3a16_PORTBDATAOUT_bus;
wire [0:0] ram_block3a49_PORTADATAOUT_bus;
wire [0:0] ram_block3a49_PORTBDATAOUT_bus;
wire [0:0] ram_block3a17_PORTADATAOUT_bus;
wire [0:0] ram_block3a17_PORTBDATAOUT_bus;
wire [0:0] ram_block3a50_PORTADATAOUT_bus;
wire [0:0] ram_block3a50_PORTBDATAOUT_bus;
wire [0:0] ram_block3a18_PORTADATAOUT_bus;
wire [0:0] ram_block3a18_PORTBDATAOUT_bus;
wire [0:0] ram_block3a51_PORTADATAOUT_bus;
wire [0:0] ram_block3a51_PORTBDATAOUT_bus;
wire [0:0] ram_block3a19_PORTADATAOUT_bus;
wire [0:0] ram_block3a19_PORTBDATAOUT_bus;
wire [0:0] ram_block3a52_PORTADATAOUT_bus;
wire [0:0] ram_block3a52_PORTBDATAOUT_bus;
wire [0:0] ram_block3a20_PORTADATAOUT_bus;
wire [0:0] ram_block3a20_PORTBDATAOUT_bus;
wire [0:0] ram_block3a53_PORTADATAOUT_bus;
wire [0:0] ram_block3a53_PORTBDATAOUT_bus;
wire [0:0] ram_block3a21_PORTADATAOUT_bus;
wire [0:0] ram_block3a21_PORTBDATAOUT_bus;
wire [0:0] ram_block3a54_PORTADATAOUT_bus;
wire [0:0] ram_block3a54_PORTBDATAOUT_bus;
wire [0:0] ram_block3a22_PORTADATAOUT_bus;
wire [0:0] ram_block3a22_PORTBDATAOUT_bus;
wire [0:0] ram_block3a55_PORTADATAOUT_bus;
wire [0:0] ram_block3a55_PORTBDATAOUT_bus;
wire [0:0] ram_block3a23_PORTADATAOUT_bus;
wire [0:0] ram_block3a23_PORTBDATAOUT_bus;
wire [0:0] ram_block3a56_PORTADATAOUT_bus;
wire [0:0] ram_block3a56_PORTBDATAOUT_bus;
wire [0:0] ram_block3a24_PORTADATAOUT_bus;
wire [0:0] ram_block3a24_PORTBDATAOUT_bus;
wire [0:0] ram_block3a57_PORTADATAOUT_bus;
wire [0:0] ram_block3a57_PORTBDATAOUT_bus;
wire [0:0] ram_block3a25_PORTADATAOUT_bus;
wire [0:0] ram_block3a25_PORTBDATAOUT_bus;
wire [0:0] ram_block3a58_PORTADATAOUT_bus;
wire [0:0] ram_block3a58_PORTBDATAOUT_bus;
wire [0:0] ram_block3a26_PORTADATAOUT_bus;
wire [0:0] ram_block3a26_PORTBDATAOUT_bus;
wire [0:0] ram_block3a59_PORTADATAOUT_bus;
wire [0:0] ram_block3a59_PORTBDATAOUT_bus;
wire [0:0] ram_block3a27_PORTADATAOUT_bus;
wire [0:0] ram_block3a27_PORTBDATAOUT_bus;
wire [0:0] ram_block3a60_PORTADATAOUT_bus;
wire [0:0] ram_block3a60_PORTBDATAOUT_bus;
wire [0:0] ram_block3a28_PORTADATAOUT_bus;
wire [0:0] ram_block3a28_PORTBDATAOUT_bus;
wire [0:0] ram_block3a61_PORTADATAOUT_bus;
wire [0:0] ram_block3a61_PORTBDATAOUT_bus;
wire [0:0] ram_block3a29_PORTADATAOUT_bus;
wire [0:0] ram_block3a29_PORTBDATAOUT_bus;
wire [0:0] ram_block3a62_PORTADATAOUT_bus;
wire [0:0] ram_block3a62_PORTBDATAOUT_bus;
wire [0:0] ram_block3a30_PORTADATAOUT_bus;
wire [0:0] ram_block3a30_PORTBDATAOUT_bus;
wire [0:0] ram_block3a63_PORTADATAOUT_bus;
wire [0:0] ram_block3a63_PORTBDATAOUT_bus;
wire [0:0] ram_block3a31_PORTADATAOUT_bus;
wire [0:0] ram_block3a31_PORTBDATAOUT_bus;

assign ram_block3a321 = ram_block3a32_PORTADATAOUT_bus[0];

assign ram_block3a322 = ram_block3a32_PORTBDATAOUT_bus[0];

assign ram_block3a01 = ram_block3a0_PORTADATAOUT_bus[0];

assign ram_block3a02 = ram_block3a0_PORTBDATAOUT_bus[0];

assign ram_block3a331 = ram_block3a33_PORTADATAOUT_bus[0];

assign ram_block3a332 = ram_block3a33_PORTBDATAOUT_bus[0];

assign ram_block3a110 = ram_block3a1_PORTADATAOUT_bus[0];

assign ram_block3a111 = ram_block3a1_PORTBDATAOUT_bus[0];

assign ram_block3a341 = ram_block3a34_PORTADATAOUT_bus[0];

assign ram_block3a342 = ram_block3a34_PORTBDATAOUT_bus[0];

assign ram_block3a210 = ram_block3a2_PORTADATAOUT_bus[0];

assign ram_block3a211 = ram_block3a2_PORTBDATAOUT_bus[0];

assign ram_block3a351 = ram_block3a35_PORTADATAOUT_bus[0];

assign ram_block3a352 = ram_block3a35_PORTBDATAOUT_bus[0];

assign ram_block3a310 = ram_block3a3_PORTADATAOUT_bus[0];

assign ram_block3a311 = ram_block3a3_PORTBDATAOUT_bus[0];

assign ram_block3a361 = ram_block3a36_PORTADATAOUT_bus[0];

assign ram_block3a362 = ram_block3a36_PORTBDATAOUT_bus[0];

assign ram_block3a410 = ram_block3a4_PORTADATAOUT_bus[0];

assign ram_block3a411 = ram_block3a4_PORTBDATAOUT_bus[0];

assign ram_block3a371 = ram_block3a37_PORTADATAOUT_bus[0];

assign ram_block3a372 = ram_block3a37_PORTBDATAOUT_bus[0];

assign ram_block3a510 = ram_block3a5_PORTADATAOUT_bus[0];

assign ram_block3a511 = ram_block3a5_PORTBDATAOUT_bus[0];

assign ram_block3a381 = ram_block3a38_PORTADATAOUT_bus[0];

assign ram_block3a382 = ram_block3a38_PORTBDATAOUT_bus[0];

assign ram_block3a64 = ram_block3a6_PORTADATAOUT_bus[0];

assign ram_block3a65 = ram_block3a6_PORTBDATAOUT_bus[0];

assign ram_block3a391 = ram_block3a39_PORTADATAOUT_bus[0];

assign ram_block3a392 = ram_block3a39_PORTBDATAOUT_bus[0];

assign ram_block3a71 = ram_block3a7_PORTADATAOUT_bus[0];

assign ram_block3a72 = ram_block3a7_PORTBDATAOUT_bus[0];

assign ram_block3a401 = ram_block3a40_PORTADATAOUT_bus[0];

assign ram_block3a402 = ram_block3a40_PORTBDATAOUT_bus[0];

assign ram_block3a81 = ram_block3a8_PORTADATAOUT_bus[0];

assign ram_block3a82 = ram_block3a8_PORTBDATAOUT_bus[0];

assign ram_block3a412 = ram_block3a41_PORTADATAOUT_bus[0];

assign ram_block3a413 = ram_block3a41_PORTBDATAOUT_bus[0];

assign ram_block3a91 = ram_block3a9_PORTADATAOUT_bus[0];

assign ram_block3a92 = ram_block3a9_PORTBDATAOUT_bus[0];

assign ram_block3a421 = ram_block3a42_PORTADATAOUT_bus[0];

assign ram_block3a422 = ram_block3a42_PORTBDATAOUT_bus[0];

assign ram_block3a101 = ram_block3a10_PORTADATAOUT_bus[0];

assign ram_block3a102 = ram_block3a10_PORTBDATAOUT_bus[0];

assign ram_block3a431 = ram_block3a43_PORTADATAOUT_bus[0];

assign ram_block3a432 = ram_block3a43_PORTBDATAOUT_bus[0];

assign ram_block3a112 = ram_block3a11_PORTADATAOUT_bus[0];

assign ram_block3a113 = ram_block3a11_PORTBDATAOUT_bus[0];

assign ram_block3a441 = ram_block3a44_PORTADATAOUT_bus[0];

assign ram_block3a442 = ram_block3a44_PORTBDATAOUT_bus[0];

assign ram_block3a121 = ram_block3a12_PORTADATAOUT_bus[0];

assign ram_block3a122 = ram_block3a12_PORTBDATAOUT_bus[0];

assign ram_block3a451 = ram_block3a45_PORTADATAOUT_bus[0];

assign ram_block3a452 = ram_block3a45_PORTBDATAOUT_bus[0];

assign ram_block3a131 = ram_block3a13_PORTADATAOUT_bus[0];

assign ram_block3a132 = ram_block3a13_PORTBDATAOUT_bus[0];

assign ram_block3a461 = ram_block3a46_PORTADATAOUT_bus[0];

assign ram_block3a462 = ram_block3a46_PORTBDATAOUT_bus[0];

assign ram_block3a141 = ram_block3a14_PORTADATAOUT_bus[0];

assign ram_block3a142 = ram_block3a14_PORTBDATAOUT_bus[0];

assign ram_block3a471 = ram_block3a47_PORTADATAOUT_bus[0];

assign ram_block3a472 = ram_block3a47_PORTBDATAOUT_bus[0];

assign ram_block3a151 = ram_block3a15_PORTADATAOUT_bus[0];

assign ram_block3a152 = ram_block3a15_PORTBDATAOUT_bus[0];

assign ram_block3a481 = ram_block3a48_PORTADATAOUT_bus[0];

assign ram_block3a482 = ram_block3a48_PORTBDATAOUT_bus[0];

assign ram_block3a161 = ram_block3a16_PORTADATAOUT_bus[0];

assign ram_block3a162 = ram_block3a16_PORTBDATAOUT_bus[0];

assign ram_block3a491 = ram_block3a49_PORTADATAOUT_bus[0];

assign ram_block3a492 = ram_block3a49_PORTBDATAOUT_bus[0];

assign ram_block3a171 = ram_block3a17_PORTADATAOUT_bus[0];

assign ram_block3a172 = ram_block3a17_PORTBDATAOUT_bus[0];

assign ram_block3a501 = ram_block3a50_PORTADATAOUT_bus[0];

assign ram_block3a502 = ram_block3a50_PORTBDATAOUT_bus[0];

assign ram_block3a181 = ram_block3a18_PORTADATAOUT_bus[0];

assign ram_block3a182 = ram_block3a18_PORTBDATAOUT_bus[0];

assign ram_block3a512 = ram_block3a51_PORTADATAOUT_bus[0];

assign ram_block3a513 = ram_block3a51_PORTBDATAOUT_bus[0];

assign ram_block3a191 = ram_block3a19_PORTADATAOUT_bus[0];

assign ram_block3a192 = ram_block3a19_PORTBDATAOUT_bus[0];

assign ram_block3a521 = ram_block3a52_PORTADATAOUT_bus[0];

assign ram_block3a522 = ram_block3a52_PORTBDATAOUT_bus[0];

assign ram_block3a201 = ram_block3a20_PORTADATAOUT_bus[0];

assign ram_block3a202 = ram_block3a20_PORTBDATAOUT_bus[0];

assign ram_block3a531 = ram_block3a53_PORTADATAOUT_bus[0];

assign ram_block3a532 = ram_block3a53_PORTBDATAOUT_bus[0];

assign ram_block3a212 = ram_block3a21_PORTADATAOUT_bus[0];

assign ram_block3a213 = ram_block3a21_PORTBDATAOUT_bus[0];

assign ram_block3a541 = ram_block3a54_PORTADATAOUT_bus[0];

assign ram_block3a542 = ram_block3a54_PORTBDATAOUT_bus[0];

assign ram_block3a221 = ram_block3a22_PORTADATAOUT_bus[0];

assign ram_block3a222 = ram_block3a22_PORTBDATAOUT_bus[0];

assign ram_block3a551 = ram_block3a55_PORTADATAOUT_bus[0];

assign ram_block3a552 = ram_block3a55_PORTBDATAOUT_bus[0];

assign ram_block3a231 = ram_block3a23_PORTADATAOUT_bus[0];

assign ram_block3a232 = ram_block3a23_PORTBDATAOUT_bus[0];

assign ram_block3a561 = ram_block3a56_PORTADATAOUT_bus[0];

assign ram_block3a562 = ram_block3a56_PORTBDATAOUT_bus[0];

assign ram_block3a241 = ram_block3a24_PORTADATAOUT_bus[0];

assign ram_block3a242 = ram_block3a24_PORTBDATAOUT_bus[0];

assign ram_block3a571 = ram_block3a57_PORTADATAOUT_bus[0];

assign ram_block3a572 = ram_block3a57_PORTBDATAOUT_bus[0];

assign ram_block3a251 = ram_block3a25_PORTADATAOUT_bus[0];

assign ram_block3a252 = ram_block3a25_PORTBDATAOUT_bus[0];

assign ram_block3a581 = ram_block3a58_PORTADATAOUT_bus[0];

assign ram_block3a582 = ram_block3a58_PORTBDATAOUT_bus[0];

assign ram_block3a261 = ram_block3a26_PORTADATAOUT_bus[0];

assign ram_block3a262 = ram_block3a26_PORTBDATAOUT_bus[0];

assign ram_block3a591 = ram_block3a59_PORTADATAOUT_bus[0];

assign ram_block3a592 = ram_block3a59_PORTBDATAOUT_bus[0];

assign ram_block3a271 = ram_block3a27_PORTADATAOUT_bus[0];

assign ram_block3a272 = ram_block3a27_PORTBDATAOUT_bus[0];

assign ram_block3a601 = ram_block3a60_PORTADATAOUT_bus[0];

assign ram_block3a602 = ram_block3a60_PORTBDATAOUT_bus[0];

assign ram_block3a281 = ram_block3a28_PORTADATAOUT_bus[0];

assign ram_block3a282 = ram_block3a28_PORTBDATAOUT_bus[0];

assign ram_block3a611 = ram_block3a61_PORTADATAOUT_bus[0];

assign ram_block3a612 = ram_block3a61_PORTBDATAOUT_bus[0];

assign ram_block3a291 = ram_block3a29_PORTADATAOUT_bus[0];

assign ram_block3a292 = ram_block3a29_PORTBDATAOUT_bus[0];

assign ram_block3a621 = ram_block3a62_PORTADATAOUT_bus[0];

assign ram_block3a622 = ram_block3a62_PORTBDATAOUT_bus[0];

assign ram_block3a301 = ram_block3a30_PORTADATAOUT_bus[0];

assign ram_block3a302 = ram_block3a30_PORTBDATAOUT_bus[0];

assign ram_block3a631 = ram_block3a63_PORTADATAOUT_bus[0];

assign ram_block3a632 = ram_block3a63_PORTBDATAOUT_bus[0];

assign ram_block3a312 = ram_block3a31_PORTADATAOUT_bus[0];

assign ram_block3a313 = ram_block3a31_PORTBDATAOUT_bus[0];

decode_jsa_1 decode5(
	.ram_rom_addr_reg_13(ram_rom_addr_reg_13),
	.sdr(sdr),
	.eq_node_1(\decode5|eq_node[1]~0_combout ),
	.eq_node_0(\decode5|eq_node[0]~1_combout ),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

decode_jsa decode4(
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.eq_node_1(\decode4|eq_node[1]~0_combout ),
	.eq_node_0(\decode4|eq_node[0]~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: M9K_X64_Y41_N0
cycloneive_ram_block ram_block3a32(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a32_PORTADATAOUT_bus),
	.portbdataout(ram_block3a32_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a32.clk0_core_clock_enable = "ena0";
defparam ram_block3a32.clk1_core_clock_enable = "ena1";
defparam ram_block3a32.data_interleave_offset_in_bits = 1;
defparam ram_block3a32.data_interleave_width_in_bits = 1;
defparam ram_block3a32.init_file = "meminit.hex";
defparam ram_block3a32.init_file_layout = "port_a";
defparam ram_block3a32.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a32.operation_mode = "bidir_dual_port";
defparam ram_block3a32.port_a_address_clear = "none";
defparam ram_block3a32.port_a_address_width = 13;
defparam ram_block3a32.port_a_byte_enable_clock = "none";
defparam ram_block3a32.port_a_data_out_clear = "none";
defparam ram_block3a32.port_a_data_out_clock = "none";
defparam ram_block3a32.port_a_data_width = 1;
defparam ram_block3a32.port_a_first_address = 0;
defparam ram_block3a32.port_a_first_bit_number = 0;
defparam ram_block3a32.port_a_last_address = 8191;
defparam ram_block3a32.port_a_logical_ram_depth = 16384;
defparam ram_block3a32.port_a_logical_ram_width = 32;
defparam ram_block3a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_address_clear = "none";
defparam ram_block3a32.port_b_address_clock = "clock1";
defparam ram_block3a32.port_b_address_width = 13;
defparam ram_block3a32.port_b_data_in_clock = "clock1";
defparam ram_block3a32.port_b_data_out_clear = "none";
defparam ram_block3a32.port_b_data_out_clock = "none";
defparam ram_block3a32.port_b_data_width = 1;
defparam ram_block3a32.port_b_first_address = 0;
defparam ram_block3a32.port_b_first_bit_number = 0;
defparam ram_block3a32.port_b_last_address = 8191;
defparam ram_block3a32.port_b_logical_ram_depth = 16384;
defparam ram_block3a32.port_b_logical_ram_width = 32;
defparam ram_block3a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_read_enable_clock = "clock1";
defparam ram_block3a32.port_b_write_enable_clock = "clock1";
defparam ram_block3a32.ram_block_type = "M9K";
defparam ram_block3a32.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y44_N0
cycloneive_ram_block ram_block3a0(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a0_PORTADATAOUT_bus),
	.portbdataout(ram_block3a0_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a0.clk0_core_clock_enable = "ena0";
defparam ram_block3a0.clk1_core_clock_enable = "ena1";
defparam ram_block3a0.data_interleave_offset_in_bits = 1;
defparam ram_block3a0.data_interleave_width_in_bits = 1;
defparam ram_block3a0.init_file = "meminit.hex";
defparam ram_block3a0.init_file_layout = "port_a";
defparam ram_block3a0.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a0.operation_mode = "bidir_dual_port";
defparam ram_block3a0.port_a_address_clear = "none";
defparam ram_block3a0.port_a_address_width = 13;
defparam ram_block3a0.port_a_byte_enable_clock = "none";
defparam ram_block3a0.port_a_data_out_clear = "none";
defparam ram_block3a0.port_a_data_out_clock = "none";
defparam ram_block3a0.port_a_data_width = 1;
defparam ram_block3a0.port_a_first_address = 0;
defparam ram_block3a0.port_a_first_bit_number = 0;
defparam ram_block3a0.port_a_last_address = 8191;
defparam ram_block3a0.port_a_logical_ram_depth = 16384;
defparam ram_block3a0.port_a_logical_ram_width = 32;
defparam ram_block3a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_address_clear = "none";
defparam ram_block3a0.port_b_address_clock = "clock1";
defparam ram_block3a0.port_b_address_width = 13;
defparam ram_block3a0.port_b_data_in_clock = "clock1";
defparam ram_block3a0.port_b_data_out_clear = "none";
defparam ram_block3a0.port_b_data_out_clock = "none";
defparam ram_block3a0.port_b_data_width = 1;
defparam ram_block3a0.port_b_first_address = 0;
defparam ram_block3a0.port_b_first_bit_number = 0;
defparam ram_block3a0.port_b_last_address = 8191;
defparam ram_block3a0.port_b_logical_ram_depth = 16384;
defparam ram_block3a0.port_b_logical_ram_width = 32;
defparam ram_block3a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_read_enable_clock = "clock1";
defparam ram_block3a0.port_b_write_enable_clock = "clock1";
defparam ram_block3a0.ram_block_type = "M9K";
defparam ram_block3a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001802C7EA14A7EF95C00000000000000000000000000000A242111E008528F7260;
// synopsys translate_on

// Location: M9K_X37_Y33_N0
cycloneive_ram_block ram_block3a33(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a33_PORTADATAOUT_bus),
	.portbdataout(ram_block3a33_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a33.clk0_core_clock_enable = "ena0";
defparam ram_block3a33.clk1_core_clock_enable = "ena1";
defparam ram_block3a33.data_interleave_offset_in_bits = 1;
defparam ram_block3a33.data_interleave_width_in_bits = 1;
defparam ram_block3a33.init_file = "meminit.hex";
defparam ram_block3a33.init_file_layout = "port_a";
defparam ram_block3a33.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a33.operation_mode = "bidir_dual_port";
defparam ram_block3a33.port_a_address_clear = "none";
defparam ram_block3a33.port_a_address_width = 13;
defparam ram_block3a33.port_a_byte_enable_clock = "none";
defparam ram_block3a33.port_a_data_out_clear = "none";
defparam ram_block3a33.port_a_data_out_clock = "none";
defparam ram_block3a33.port_a_data_width = 1;
defparam ram_block3a33.port_a_first_address = 0;
defparam ram_block3a33.port_a_first_bit_number = 1;
defparam ram_block3a33.port_a_last_address = 8191;
defparam ram_block3a33.port_a_logical_ram_depth = 16384;
defparam ram_block3a33.port_a_logical_ram_width = 32;
defparam ram_block3a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_address_clear = "none";
defparam ram_block3a33.port_b_address_clock = "clock1";
defparam ram_block3a33.port_b_address_width = 13;
defparam ram_block3a33.port_b_data_in_clock = "clock1";
defparam ram_block3a33.port_b_data_out_clear = "none";
defparam ram_block3a33.port_b_data_out_clock = "none";
defparam ram_block3a33.port_b_data_width = 1;
defparam ram_block3a33.port_b_first_address = 0;
defparam ram_block3a33.port_b_first_bit_number = 1;
defparam ram_block3a33.port_b_last_address = 8191;
defparam ram_block3a33.port_b_logical_ram_depth = 16384;
defparam ram_block3a33.port_b_logical_ram_width = 32;
defparam ram_block3a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_read_enable_clock = "clock1";
defparam ram_block3a33.port_b_write_enable_clock = "clock1";
defparam ram_block3a33.ram_block_type = "M9K";
defparam ram_block3a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y36_N0
cycloneive_ram_block ram_block3a1(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a1_PORTADATAOUT_bus),
	.portbdataout(ram_block3a1_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a1.clk0_core_clock_enable = "ena0";
defparam ram_block3a1.clk1_core_clock_enable = "ena1";
defparam ram_block3a1.data_interleave_offset_in_bits = 1;
defparam ram_block3a1.data_interleave_width_in_bits = 1;
defparam ram_block3a1.init_file = "meminit.hex";
defparam ram_block3a1.init_file_layout = "port_a";
defparam ram_block3a1.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a1.operation_mode = "bidir_dual_port";
defparam ram_block3a1.port_a_address_clear = "none";
defparam ram_block3a1.port_a_address_width = 13;
defparam ram_block3a1.port_a_byte_enable_clock = "none";
defparam ram_block3a1.port_a_data_out_clear = "none";
defparam ram_block3a1.port_a_data_out_clock = "none";
defparam ram_block3a1.port_a_data_width = 1;
defparam ram_block3a1.port_a_first_address = 0;
defparam ram_block3a1.port_a_first_bit_number = 1;
defparam ram_block3a1.port_a_last_address = 8191;
defparam ram_block3a1.port_a_logical_ram_depth = 16384;
defparam ram_block3a1.port_a_logical_ram_width = 32;
defparam ram_block3a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_address_clear = "none";
defparam ram_block3a1.port_b_address_clock = "clock1";
defparam ram_block3a1.port_b_address_width = 13;
defparam ram_block3a1.port_b_data_in_clock = "clock1";
defparam ram_block3a1.port_b_data_out_clear = "none";
defparam ram_block3a1.port_b_data_out_clock = "none";
defparam ram_block3a1.port_b_data_width = 1;
defparam ram_block3a1.port_b_first_address = 0;
defparam ram_block3a1.port_b_first_bit_number = 1;
defparam ram_block3a1.port_b_last_address = 8191;
defparam ram_block3a1.port_b_logical_ram_depth = 16384;
defparam ram_block3a1.port_b_logical_ram_width = 32;
defparam ram_block3a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_read_enable_clock = "clock1";
defparam ram_block3a1.port_b_write_enable_clock = "clock1";
defparam ram_block3a1.ram_block_type = "M9K";
defparam ram_block3a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001D4AE6429116B3C8A000000000000000000000000000012242108900D12808390;
// synopsys translate_on

// Location: M9K_X37_Y35_N0
cycloneive_ram_block ram_block3a34(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a34_PORTADATAOUT_bus),
	.portbdataout(ram_block3a34_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a34.clk0_core_clock_enable = "ena0";
defparam ram_block3a34.clk1_core_clock_enable = "ena1";
defparam ram_block3a34.data_interleave_offset_in_bits = 1;
defparam ram_block3a34.data_interleave_width_in_bits = 1;
defparam ram_block3a34.init_file = "meminit.hex";
defparam ram_block3a34.init_file_layout = "port_a";
defparam ram_block3a34.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a34.operation_mode = "bidir_dual_port";
defparam ram_block3a34.port_a_address_clear = "none";
defparam ram_block3a34.port_a_address_width = 13;
defparam ram_block3a34.port_a_byte_enable_clock = "none";
defparam ram_block3a34.port_a_data_out_clear = "none";
defparam ram_block3a34.port_a_data_out_clock = "none";
defparam ram_block3a34.port_a_data_width = 1;
defparam ram_block3a34.port_a_first_address = 0;
defparam ram_block3a34.port_a_first_bit_number = 2;
defparam ram_block3a34.port_a_last_address = 8191;
defparam ram_block3a34.port_a_logical_ram_depth = 16384;
defparam ram_block3a34.port_a_logical_ram_width = 32;
defparam ram_block3a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_address_clear = "none";
defparam ram_block3a34.port_b_address_clock = "clock1";
defparam ram_block3a34.port_b_address_width = 13;
defparam ram_block3a34.port_b_data_in_clock = "clock1";
defparam ram_block3a34.port_b_data_out_clear = "none";
defparam ram_block3a34.port_b_data_out_clock = "none";
defparam ram_block3a34.port_b_data_width = 1;
defparam ram_block3a34.port_b_first_address = 0;
defparam ram_block3a34.port_b_first_bit_number = 2;
defparam ram_block3a34.port_b_last_address = 8191;
defparam ram_block3a34.port_b_logical_ram_depth = 16384;
defparam ram_block3a34.port_b_logical_ram_width = 32;
defparam ram_block3a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_read_enable_clock = "clock1";
defparam ram_block3a34.port_b_write_enable_clock = "clock1";
defparam ram_block3a34.ram_block_type = "M9K";
defparam ram_block3a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y30_N0
cycloneive_ram_block ram_block3a2(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a2_PORTADATAOUT_bus),
	.portbdataout(ram_block3a2_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a2.clk0_core_clock_enable = "ena0";
defparam ram_block3a2.clk1_core_clock_enable = "ena1";
defparam ram_block3a2.data_interleave_offset_in_bits = 1;
defparam ram_block3a2.data_interleave_width_in_bits = 1;
defparam ram_block3a2.init_file = "meminit.hex";
defparam ram_block3a2.init_file_layout = "port_a";
defparam ram_block3a2.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a2.operation_mode = "bidir_dual_port";
defparam ram_block3a2.port_a_address_clear = "none";
defparam ram_block3a2.port_a_address_width = 13;
defparam ram_block3a2.port_a_byte_enable_clock = "none";
defparam ram_block3a2.port_a_data_out_clear = "none";
defparam ram_block3a2.port_a_data_out_clock = "none";
defparam ram_block3a2.port_a_data_width = 1;
defparam ram_block3a2.port_a_first_address = 0;
defparam ram_block3a2.port_a_first_bit_number = 2;
defparam ram_block3a2.port_a_last_address = 8191;
defparam ram_block3a2.port_a_logical_ram_depth = 16384;
defparam ram_block3a2.port_a_logical_ram_width = 32;
defparam ram_block3a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_address_clear = "none";
defparam ram_block3a2.port_b_address_clock = "clock1";
defparam ram_block3a2.port_b_address_width = 13;
defparam ram_block3a2.port_b_data_in_clock = "clock1";
defparam ram_block3a2.port_b_data_out_clear = "none";
defparam ram_block3a2.port_b_data_out_clock = "none";
defparam ram_block3a2.port_b_data_width = 1;
defparam ram_block3a2.port_b_first_address = 0;
defparam ram_block3a2.port_b_first_bit_number = 2;
defparam ram_block3a2.port_b_last_address = 8191;
defparam ram_block3a2.port_b_logical_ram_depth = 16384;
defparam ram_block3a2.port_b_logical_ram_width = 32;
defparam ram_block3a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_read_enable_clock = "clock1";
defparam ram_block3a2.port_b_write_enable_clock = "clock1";
defparam ram_block3a2.ram_block_type = "M9K";
defparam ram_block3a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000961CA470728D97800000000000000000000000000000172E7BD1C323272F6867;
// synopsys translate_on

// Location: M9K_X64_Y43_N0
cycloneive_ram_block ram_block3a35(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a35_PORTADATAOUT_bus),
	.portbdataout(ram_block3a35_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a35.clk0_core_clock_enable = "ena0";
defparam ram_block3a35.clk1_core_clock_enable = "ena1";
defparam ram_block3a35.data_interleave_offset_in_bits = 1;
defparam ram_block3a35.data_interleave_width_in_bits = 1;
defparam ram_block3a35.init_file = "meminit.hex";
defparam ram_block3a35.init_file_layout = "port_a";
defparam ram_block3a35.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a35.operation_mode = "bidir_dual_port";
defparam ram_block3a35.port_a_address_clear = "none";
defparam ram_block3a35.port_a_address_width = 13;
defparam ram_block3a35.port_a_byte_enable_clock = "none";
defparam ram_block3a35.port_a_data_out_clear = "none";
defparam ram_block3a35.port_a_data_out_clock = "none";
defparam ram_block3a35.port_a_data_width = 1;
defparam ram_block3a35.port_a_first_address = 0;
defparam ram_block3a35.port_a_first_bit_number = 3;
defparam ram_block3a35.port_a_last_address = 8191;
defparam ram_block3a35.port_a_logical_ram_depth = 16384;
defparam ram_block3a35.port_a_logical_ram_width = 32;
defparam ram_block3a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_address_clear = "none";
defparam ram_block3a35.port_b_address_clock = "clock1";
defparam ram_block3a35.port_b_address_width = 13;
defparam ram_block3a35.port_b_data_in_clock = "clock1";
defparam ram_block3a35.port_b_data_out_clear = "none";
defparam ram_block3a35.port_b_data_out_clock = "none";
defparam ram_block3a35.port_b_data_width = 1;
defparam ram_block3a35.port_b_first_address = 0;
defparam ram_block3a35.port_b_first_bit_number = 3;
defparam ram_block3a35.port_b_last_address = 8191;
defparam ram_block3a35.port_b_logical_ram_depth = 16384;
defparam ram_block3a35.port_b_logical_ram_width = 32;
defparam ram_block3a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_read_enable_clock = "clock1";
defparam ram_block3a35.port_b_write_enable_clock = "clock1";
defparam ram_block3a35.ram_block_type = "M9K";
defparam ram_block3a35.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y46_N0
cycloneive_ram_block ram_block3a3(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a3_PORTADATAOUT_bus),
	.portbdataout(ram_block3a3_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a3.clk0_core_clock_enable = "ena0";
defparam ram_block3a3.clk1_core_clock_enable = "ena1";
defparam ram_block3a3.data_interleave_offset_in_bits = 1;
defparam ram_block3a3.data_interleave_width_in_bits = 1;
defparam ram_block3a3.init_file = "meminit.hex";
defparam ram_block3a3.init_file_layout = "port_a";
defparam ram_block3a3.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a3.operation_mode = "bidir_dual_port";
defparam ram_block3a3.port_a_address_clear = "none";
defparam ram_block3a3.port_a_address_width = 13;
defparam ram_block3a3.port_a_byte_enable_clock = "none";
defparam ram_block3a3.port_a_data_out_clear = "none";
defparam ram_block3a3.port_a_data_out_clock = "none";
defparam ram_block3a3.port_a_data_width = 1;
defparam ram_block3a3.port_a_first_address = 0;
defparam ram_block3a3.port_a_first_bit_number = 3;
defparam ram_block3a3.port_a_last_address = 8191;
defparam ram_block3a3.port_a_logical_ram_depth = 16384;
defparam ram_block3a3.port_a_logical_ram_width = 32;
defparam ram_block3a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_address_clear = "none";
defparam ram_block3a3.port_b_address_clock = "clock1";
defparam ram_block3a3.port_b_address_width = 13;
defparam ram_block3a3.port_b_data_in_clock = "clock1";
defparam ram_block3a3.port_b_data_out_clear = "none";
defparam ram_block3a3.port_b_data_out_clock = "none";
defparam ram_block3a3.port_b_data_width = 1;
defparam ram_block3a3.port_b_first_address = 0;
defparam ram_block3a3.port_b_first_bit_number = 3;
defparam ram_block3a3.port_b_last_address = 8191;
defparam ram_block3a3.port_b_logical_ram_depth = 16384;
defparam ram_block3a3.port_b_logical_ram_width = 32;
defparam ram_block3a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_read_enable_clock = "clock1";
defparam ram_block3a3.port_b_write_enable_clock = "clock1";
defparam ram_block3a3.ram_block_type = "M9K";
defparam ram_block3a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009F20E64C2468E52000000000000000000000000000022346308C62632A08083;
// synopsys translate_on

// Location: M9K_X64_Y48_N0
cycloneive_ram_block ram_block3a36(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a36_PORTADATAOUT_bus),
	.portbdataout(ram_block3a36_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a36.clk0_core_clock_enable = "ena0";
defparam ram_block3a36.clk1_core_clock_enable = "ena1";
defparam ram_block3a36.data_interleave_offset_in_bits = 1;
defparam ram_block3a36.data_interleave_width_in_bits = 1;
defparam ram_block3a36.init_file = "meminit.hex";
defparam ram_block3a36.init_file_layout = "port_a";
defparam ram_block3a36.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a36.operation_mode = "bidir_dual_port";
defparam ram_block3a36.port_a_address_clear = "none";
defparam ram_block3a36.port_a_address_width = 13;
defparam ram_block3a36.port_a_byte_enable_clock = "none";
defparam ram_block3a36.port_a_data_out_clear = "none";
defparam ram_block3a36.port_a_data_out_clock = "none";
defparam ram_block3a36.port_a_data_width = 1;
defparam ram_block3a36.port_a_first_address = 0;
defparam ram_block3a36.port_a_first_bit_number = 4;
defparam ram_block3a36.port_a_last_address = 8191;
defparam ram_block3a36.port_a_logical_ram_depth = 16384;
defparam ram_block3a36.port_a_logical_ram_width = 32;
defparam ram_block3a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_address_clear = "none";
defparam ram_block3a36.port_b_address_clock = "clock1";
defparam ram_block3a36.port_b_address_width = 13;
defparam ram_block3a36.port_b_data_in_clock = "clock1";
defparam ram_block3a36.port_b_data_out_clear = "none";
defparam ram_block3a36.port_b_data_out_clock = "none";
defparam ram_block3a36.port_b_data_width = 1;
defparam ram_block3a36.port_b_first_address = 0;
defparam ram_block3a36.port_b_first_bit_number = 4;
defparam ram_block3a36.port_b_last_address = 8191;
defparam ram_block3a36.port_b_logical_ram_depth = 16384;
defparam ram_block3a36.port_b_logical_ram_width = 32;
defparam ram_block3a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_read_enable_clock = "clock1";
defparam ram_block3a36.port_b_write_enable_clock = "clock1";
defparam ram_block3a36.ram_block_type = "M9K";
defparam ram_block3a36.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y47_N0
cycloneive_ram_block ram_block3a4(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a4_PORTADATAOUT_bus),
	.portbdataout(ram_block3a4_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a4.clk0_core_clock_enable = "ena0";
defparam ram_block3a4.clk1_core_clock_enable = "ena1";
defparam ram_block3a4.data_interleave_offset_in_bits = 1;
defparam ram_block3a4.data_interleave_width_in_bits = 1;
defparam ram_block3a4.init_file = "meminit.hex";
defparam ram_block3a4.init_file_layout = "port_a";
defparam ram_block3a4.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a4.operation_mode = "bidir_dual_port";
defparam ram_block3a4.port_a_address_clear = "none";
defparam ram_block3a4.port_a_address_width = 13;
defparam ram_block3a4.port_a_byte_enable_clock = "none";
defparam ram_block3a4.port_a_data_out_clear = "none";
defparam ram_block3a4.port_a_data_out_clock = "none";
defparam ram_block3a4.port_a_data_width = 1;
defparam ram_block3a4.port_a_first_address = 0;
defparam ram_block3a4.port_a_first_bit_number = 4;
defparam ram_block3a4.port_a_last_address = 8191;
defparam ram_block3a4.port_a_logical_ram_depth = 16384;
defparam ram_block3a4.port_a_logical_ram_width = 32;
defparam ram_block3a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_address_clear = "none";
defparam ram_block3a4.port_b_address_clock = "clock1";
defparam ram_block3a4.port_b_address_width = 13;
defparam ram_block3a4.port_b_data_in_clock = "clock1";
defparam ram_block3a4.port_b_data_out_clear = "none";
defparam ram_block3a4.port_b_data_out_clock = "none";
defparam ram_block3a4.port_b_data_width = 1;
defparam ram_block3a4.port_b_first_address = 0;
defparam ram_block3a4.port_b_first_bit_number = 4;
defparam ram_block3a4.port_b_last_address = 8191;
defparam ram_block3a4.port_b_logical_ram_depth = 16384;
defparam ram_block3a4.port_b_logical_ram_width = 32;
defparam ram_block3a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_read_enable_clock = "clock1";
defparam ram_block3a4.port_b_write_enable_clock = "clock1";
defparam ram_block3a4.ram_block_type = "M9K";
defparam ram_block3a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060B81842D24565BE000000000000000000000000000002242101022202208083;
// synopsys translate_on

// Location: M9K_X64_Y30_N0
cycloneive_ram_block ram_block3a37(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a37_PORTADATAOUT_bus),
	.portbdataout(ram_block3a37_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a37.clk0_core_clock_enable = "ena0";
defparam ram_block3a37.clk1_core_clock_enable = "ena1";
defparam ram_block3a37.data_interleave_offset_in_bits = 1;
defparam ram_block3a37.data_interleave_width_in_bits = 1;
defparam ram_block3a37.init_file = "meminit.hex";
defparam ram_block3a37.init_file_layout = "port_a";
defparam ram_block3a37.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a37.operation_mode = "bidir_dual_port";
defparam ram_block3a37.port_a_address_clear = "none";
defparam ram_block3a37.port_a_address_width = 13;
defparam ram_block3a37.port_a_byte_enable_clock = "none";
defparam ram_block3a37.port_a_data_out_clear = "none";
defparam ram_block3a37.port_a_data_out_clock = "none";
defparam ram_block3a37.port_a_data_width = 1;
defparam ram_block3a37.port_a_first_address = 0;
defparam ram_block3a37.port_a_first_bit_number = 5;
defparam ram_block3a37.port_a_last_address = 8191;
defparam ram_block3a37.port_a_logical_ram_depth = 16384;
defparam ram_block3a37.port_a_logical_ram_width = 32;
defparam ram_block3a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_address_clear = "none";
defparam ram_block3a37.port_b_address_clock = "clock1";
defparam ram_block3a37.port_b_address_width = 13;
defparam ram_block3a37.port_b_data_in_clock = "clock1";
defparam ram_block3a37.port_b_data_out_clear = "none";
defparam ram_block3a37.port_b_data_out_clock = "none";
defparam ram_block3a37.port_b_data_width = 1;
defparam ram_block3a37.port_b_first_address = 0;
defparam ram_block3a37.port_b_first_bit_number = 5;
defparam ram_block3a37.port_b_last_address = 8191;
defparam ram_block3a37.port_b_logical_ram_depth = 16384;
defparam ram_block3a37.port_b_logical_ram_width = 32;
defparam ram_block3a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_read_enable_clock = "clock1";
defparam ram_block3a37.port_b_write_enable_clock = "clock1";
defparam ram_block3a37.ram_block_type = "M9K";
defparam ram_block3a37.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y31_N0
cycloneive_ram_block ram_block3a5(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a5_PORTADATAOUT_bus),
	.portbdataout(ram_block3a5_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a5.clk0_core_clock_enable = "ena0";
defparam ram_block3a5.clk1_core_clock_enable = "ena1";
defparam ram_block3a5.data_interleave_offset_in_bits = 1;
defparam ram_block3a5.data_interleave_width_in_bits = 1;
defparam ram_block3a5.init_file = "meminit.hex";
defparam ram_block3a5.init_file_layout = "port_a";
defparam ram_block3a5.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a5.operation_mode = "bidir_dual_port";
defparam ram_block3a5.port_a_address_clear = "none";
defparam ram_block3a5.port_a_address_width = 13;
defparam ram_block3a5.port_a_byte_enable_clock = "none";
defparam ram_block3a5.port_a_data_out_clear = "none";
defparam ram_block3a5.port_a_data_out_clock = "none";
defparam ram_block3a5.port_a_data_width = 1;
defparam ram_block3a5.port_a_first_address = 0;
defparam ram_block3a5.port_a_first_bit_number = 5;
defparam ram_block3a5.port_a_last_address = 8191;
defparam ram_block3a5.port_a_logical_ram_depth = 16384;
defparam ram_block3a5.port_a_logical_ram_width = 32;
defparam ram_block3a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_address_clear = "none";
defparam ram_block3a5.port_b_address_clock = "clock1";
defparam ram_block3a5.port_b_address_width = 13;
defparam ram_block3a5.port_b_data_in_clock = "clock1";
defparam ram_block3a5.port_b_data_out_clear = "none";
defparam ram_block3a5.port_b_data_out_clock = "none";
defparam ram_block3a5.port_b_data_width = 1;
defparam ram_block3a5.port_b_first_address = 0;
defparam ram_block3a5.port_b_first_bit_number = 5;
defparam ram_block3a5.port_b_last_address = 8191;
defparam ram_block3a5.port_b_logical_ram_depth = 16384;
defparam ram_block3a5.port_b_logical_ram_width = 32;
defparam ram_block3a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_read_enable_clock = "clock1";
defparam ram_block3a5.port_b_write_enable_clock = "clock1";
defparam ram_block3a5.ram_block_type = "M9K";
defparam ram_block3a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000056414512D6B00448000000000000000000000000000002246308006652AF7263;
// synopsys translate_on

// Location: M9K_X78_Y32_N0
cycloneive_ram_block ram_block3a38(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a38_PORTADATAOUT_bus),
	.portbdataout(ram_block3a38_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a38.clk0_core_clock_enable = "ena0";
defparam ram_block3a38.clk1_core_clock_enable = "ena1";
defparam ram_block3a38.data_interleave_offset_in_bits = 1;
defparam ram_block3a38.data_interleave_width_in_bits = 1;
defparam ram_block3a38.init_file = "meminit.hex";
defparam ram_block3a38.init_file_layout = "port_a";
defparam ram_block3a38.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a38.operation_mode = "bidir_dual_port";
defparam ram_block3a38.port_a_address_clear = "none";
defparam ram_block3a38.port_a_address_width = 13;
defparam ram_block3a38.port_a_byte_enable_clock = "none";
defparam ram_block3a38.port_a_data_out_clear = "none";
defparam ram_block3a38.port_a_data_out_clock = "none";
defparam ram_block3a38.port_a_data_width = 1;
defparam ram_block3a38.port_a_first_address = 0;
defparam ram_block3a38.port_a_first_bit_number = 6;
defparam ram_block3a38.port_a_last_address = 8191;
defparam ram_block3a38.port_a_logical_ram_depth = 16384;
defparam ram_block3a38.port_a_logical_ram_width = 32;
defparam ram_block3a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_address_clear = "none";
defparam ram_block3a38.port_b_address_clock = "clock1";
defparam ram_block3a38.port_b_address_width = 13;
defparam ram_block3a38.port_b_data_in_clock = "clock1";
defparam ram_block3a38.port_b_data_out_clear = "none";
defparam ram_block3a38.port_b_data_out_clock = "none";
defparam ram_block3a38.port_b_data_width = 1;
defparam ram_block3a38.port_b_first_address = 0;
defparam ram_block3a38.port_b_first_bit_number = 6;
defparam ram_block3a38.port_b_last_address = 8191;
defparam ram_block3a38.port_b_logical_ram_depth = 16384;
defparam ram_block3a38.port_b_logical_ram_width = 32;
defparam ram_block3a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_read_enable_clock = "clock1";
defparam ram_block3a38.port_b_write_enable_clock = "clock1";
defparam ram_block3a38.ram_block_type = "M9K";
defparam ram_block3a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y31_N0
cycloneive_ram_block ram_block3a6(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a6_PORTADATAOUT_bus),
	.portbdataout(ram_block3a6_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a6.clk0_core_clock_enable = "ena0";
defparam ram_block3a6.clk1_core_clock_enable = "ena1";
defparam ram_block3a6.data_interleave_offset_in_bits = 1;
defparam ram_block3a6.data_interleave_width_in_bits = 1;
defparam ram_block3a6.init_file = "meminit.hex";
defparam ram_block3a6.init_file_layout = "port_a";
defparam ram_block3a6.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a6.operation_mode = "bidir_dual_port";
defparam ram_block3a6.port_a_address_clear = "none";
defparam ram_block3a6.port_a_address_width = 13;
defparam ram_block3a6.port_a_byte_enable_clock = "none";
defparam ram_block3a6.port_a_data_out_clear = "none";
defparam ram_block3a6.port_a_data_out_clock = "none";
defparam ram_block3a6.port_a_data_width = 1;
defparam ram_block3a6.port_a_first_address = 0;
defparam ram_block3a6.port_a_first_bit_number = 6;
defparam ram_block3a6.port_a_last_address = 8191;
defparam ram_block3a6.port_a_logical_ram_depth = 16384;
defparam ram_block3a6.port_a_logical_ram_width = 32;
defparam ram_block3a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_address_clear = "none";
defparam ram_block3a6.port_b_address_clock = "clock1";
defparam ram_block3a6.port_b_address_width = 13;
defparam ram_block3a6.port_b_data_in_clock = "clock1";
defparam ram_block3a6.port_b_data_out_clear = "none";
defparam ram_block3a6.port_b_data_out_clock = "none";
defparam ram_block3a6.port_b_data_width = 1;
defparam ram_block3a6.port_b_first_address = 0;
defparam ram_block3a6.port_b_first_bit_number = 6;
defparam ram_block3a6.port_b_last_address = 8191;
defparam ram_block3a6.port_b_logical_ram_depth = 16384;
defparam ram_block3a6.port_b_logical_ram_width = 32;
defparam ram_block3a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_read_enable_clock = "clock1";
defparam ram_block3a6.port_b_write_enable_clock = "clock1";
defparam ram_block3a6.ram_block_type = "M9K";
defparam ram_block3a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001003088D801A0F827000000000000000000000000000012042100402202200113;
// synopsys translate_on

// Location: M9K_X37_Y34_N0
cycloneive_ram_block ram_block3a39(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a39_PORTADATAOUT_bus),
	.portbdataout(ram_block3a39_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a39.clk0_core_clock_enable = "ena0";
defparam ram_block3a39.clk1_core_clock_enable = "ena1";
defparam ram_block3a39.data_interleave_offset_in_bits = 1;
defparam ram_block3a39.data_interleave_width_in_bits = 1;
defparam ram_block3a39.init_file = "meminit.hex";
defparam ram_block3a39.init_file_layout = "port_a";
defparam ram_block3a39.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a39.operation_mode = "bidir_dual_port";
defparam ram_block3a39.port_a_address_clear = "none";
defparam ram_block3a39.port_a_address_width = 13;
defparam ram_block3a39.port_a_byte_enable_clock = "none";
defparam ram_block3a39.port_a_data_out_clear = "none";
defparam ram_block3a39.port_a_data_out_clock = "none";
defparam ram_block3a39.port_a_data_width = 1;
defparam ram_block3a39.port_a_first_address = 0;
defparam ram_block3a39.port_a_first_bit_number = 7;
defparam ram_block3a39.port_a_last_address = 8191;
defparam ram_block3a39.port_a_logical_ram_depth = 16384;
defparam ram_block3a39.port_a_logical_ram_width = 32;
defparam ram_block3a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_address_clear = "none";
defparam ram_block3a39.port_b_address_clock = "clock1";
defparam ram_block3a39.port_b_address_width = 13;
defparam ram_block3a39.port_b_data_in_clock = "clock1";
defparam ram_block3a39.port_b_data_out_clear = "none";
defparam ram_block3a39.port_b_data_out_clock = "none";
defparam ram_block3a39.port_b_data_width = 1;
defparam ram_block3a39.port_b_first_address = 0;
defparam ram_block3a39.port_b_first_bit_number = 7;
defparam ram_block3a39.port_b_last_address = 8191;
defparam ram_block3a39.port_b_logical_ram_depth = 16384;
defparam ram_block3a39.port_b_logical_ram_width = 32;
defparam ram_block3a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_read_enable_clock = "clock1";
defparam ram_block3a39.port_b_write_enable_clock = "clock1";
defparam ram_block3a39.ram_block_type = "M9K";
defparam ram_block3a39.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y38_N0
cycloneive_ram_block ram_block3a7(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a7_PORTADATAOUT_bus),
	.portbdataout(ram_block3a7_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a7.clk0_core_clock_enable = "ena0";
defparam ram_block3a7.clk1_core_clock_enable = "ena1";
defparam ram_block3a7.data_interleave_offset_in_bits = 1;
defparam ram_block3a7.data_interleave_width_in_bits = 1;
defparam ram_block3a7.init_file = "meminit.hex";
defparam ram_block3a7.init_file_layout = "port_a";
defparam ram_block3a7.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a7.operation_mode = "bidir_dual_port";
defparam ram_block3a7.port_a_address_clear = "none";
defparam ram_block3a7.port_a_address_width = 13;
defparam ram_block3a7.port_a_byte_enable_clock = "none";
defparam ram_block3a7.port_a_data_out_clear = "none";
defparam ram_block3a7.port_a_data_out_clock = "none";
defparam ram_block3a7.port_a_data_width = 1;
defparam ram_block3a7.port_a_first_address = 0;
defparam ram_block3a7.port_a_first_bit_number = 7;
defparam ram_block3a7.port_a_last_address = 8191;
defparam ram_block3a7.port_a_logical_ram_depth = 16384;
defparam ram_block3a7.port_a_logical_ram_width = 32;
defparam ram_block3a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_address_clear = "none";
defparam ram_block3a7.port_b_address_clock = "clock1";
defparam ram_block3a7.port_b_address_width = 13;
defparam ram_block3a7.port_b_data_in_clock = "clock1";
defparam ram_block3a7.port_b_data_out_clear = "none";
defparam ram_block3a7.port_b_data_out_clock = "none";
defparam ram_block3a7.port_b_data_width = 1;
defparam ram_block3a7.port_b_first_address = 0;
defparam ram_block3a7.port_b_first_bit_number = 7;
defparam ram_block3a7.port_b_last_address = 8191;
defparam ram_block3a7.port_b_logical_ram_depth = 16384;
defparam ram_block3a7.port_b_logical_ram_width = 32;
defparam ram_block3a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_read_enable_clock = "clock1";
defparam ram_block3a7.port_b_write_enable_clock = "clock1";
defparam ram_block3a7.ram_block_type = "M9K";
defparam ram_block3a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220A200403;
// synopsys translate_on

// Location: M9K_X78_Y34_N0
cycloneive_ram_block ram_block3a40(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a40_PORTADATAOUT_bus),
	.portbdataout(ram_block3a40_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a40.clk0_core_clock_enable = "ena0";
defparam ram_block3a40.clk1_core_clock_enable = "ena1";
defparam ram_block3a40.data_interleave_offset_in_bits = 1;
defparam ram_block3a40.data_interleave_width_in_bits = 1;
defparam ram_block3a40.init_file = "meminit.hex";
defparam ram_block3a40.init_file_layout = "port_a";
defparam ram_block3a40.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a40.operation_mode = "bidir_dual_port";
defparam ram_block3a40.port_a_address_clear = "none";
defparam ram_block3a40.port_a_address_width = 13;
defparam ram_block3a40.port_a_byte_enable_clock = "none";
defparam ram_block3a40.port_a_data_out_clear = "none";
defparam ram_block3a40.port_a_data_out_clock = "none";
defparam ram_block3a40.port_a_data_width = 1;
defparam ram_block3a40.port_a_first_address = 0;
defparam ram_block3a40.port_a_first_bit_number = 8;
defparam ram_block3a40.port_a_last_address = 8191;
defparam ram_block3a40.port_a_logical_ram_depth = 16384;
defparam ram_block3a40.port_a_logical_ram_width = 32;
defparam ram_block3a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_address_clear = "none";
defparam ram_block3a40.port_b_address_clock = "clock1";
defparam ram_block3a40.port_b_address_width = 13;
defparam ram_block3a40.port_b_data_in_clock = "clock1";
defparam ram_block3a40.port_b_data_out_clear = "none";
defparam ram_block3a40.port_b_data_out_clock = "none";
defparam ram_block3a40.port_b_data_width = 1;
defparam ram_block3a40.port_b_first_address = 0;
defparam ram_block3a40.port_b_first_bit_number = 8;
defparam ram_block3a40.port_b_last_address = 8191;
defparam ram_block3a40.port_b_logical_ram_depth = 16384;
defparam ram_block3a40.port_b_logical_ram_width = 32;
defparam ram_block3a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_read_enable_clock = "clock1";
defparam ram_block3a40.port_b_write_enable_clock = "clock1";
defparam ram_block3a40.ram_block_type = "M9K";
defparam ram_block3a40.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y35_N0
cycloneive_ram_block ram_block3a8(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a8_PORTADATAOUT_bus),
	.portbdataout(ram_block3a8_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a8.clk0_core_clock_enable = "ena0";
defparam ram_block3a8.clk1_core_clock_enable = "ena1";
defparam ram_block3a8.data_interleave_offset_in_bits = 1;
defparam ram_block3a8.data_interleave_width_in_bits = 1;
defparam ram_block3a8.init_file = "meminit.hex";
defparam ram_block3a8.init_file_layout = "port_a";
defparam ram_block3a8.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a8.operation_mode = "bidir_dual_port";
defparam ram_block3a8.port_a_address_clear = "none";
defparam ram_block3a8.port_a_address_width = 13;
defparam ram_block3a8.port_a_byte_enable_clock = "none";
defparam ram_block3a8.port_a_data_out_clear = "none";
defparam ram_block3a8.port_a_data_out_clock = "none";
defparam ram_block3a8.port_a_data_width = 1;
defparam ram_block3a8.port_a_first_address = 0;
defparam ram_block3a8.port_a_first_bit_number = 8;
defparam ram_block3a8.port_a_last_address = 8191;
defparam ram_block3a8.port_a_logical_ram_depth = 16384;
defparam ram_block3a8.port_a_logical_ram_width = 32;
defparam ram_block3a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_address_clear = "none";
defparam ram_block3a8.port_b_address_clock = "clock1";
defparam ram_block3a8.port_b_address_width = 13;
defparam ram_block3a8.port_b_data_in_clock = "clock1";
defparam ram_block3a8.port_b_data_out_clear = "none";
defparam ram_block3a8.port_b_data_out_clock = "none";
defparam ram_block3a8.port_b_data_width = 1;
defparam ram_block3a8.port_b_first_address = 0;
defparam ram_block3a8.port_b_first_bit_number = 8;
defparam ram_block3a8.port_b_last_address = 8191;
defparam ram_block3a8.port_b_logical_ram_depth = 16384;
defparam ram_block3a8.port_b_logical_ram_width = 32;
defparam ram_block3a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_read_enable_clock = "clock1";
defparam ram_block3a8.port_b_write_enable_clock = "clock1";
defparam ram_block3a8.ram_block_type = "M9K";
defparam ram_block3a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220230080F;
// synopsys translate_on

// Location: M9K_X78_Y43_N0
cycloneive_ram_block ram_block3a41(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a41_PORTADATAOUT_bus),
	.portbdataout(ram_block3a41_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a41.clk0_core_clock_enable = "ena0";
defparam ram_block3a41.clk1_core_clock_enable = "ena1";
defparam ram_block3a41.data_interleave_offset_in_bits = 1;
defparam ram_block3a41.data_interleave_width_in_bits = 1;
defparam ram_block3a41.init_file = "meminit.hex";
defparam ram_block3a41.init_file_layout = "port_a";
defparam ram_block3a41.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a41.operation_mode = "bidir_dual_port";
defparam ram_block3a41.port_a_address_clear = "none";
defparam ram_block3a41.port_a_address_width = 13;
defparam ram_block3a41.port_a_byte_enable_clock = "none";
defparam ram_block3a41.port_a_data_out_clear = "none";
defparam ram_block3a41.port_a_data_out_clock = "none";
defparam ram_block3a41.port_a_data_width = 1;
defparam ram_block3a41.port_a_first_address = 0;
defparam ram_block3a41.port_a_first_bit_number = 9;
defparam ram_block3a41.port_a_last_address = 8191;
defparam ram_block3a41.port_a_logical_ram_depth = 16384;
defparam ram_block3a41.port_a_logical_ram_width = 32;
defparam ram_block3a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_address_clear = "none";
defparam ram_block3a41.port_b_address_clock = "clock1";
defparam ram_block3a41.port_b_address_width = 13;
defparam ram_block3a41.port_b_data_in_clock = "clock1";
defparam ram_block3a41.port_b_data_out_clear = "none";
defparam ram_block3a41.port_b_data_out_clock = "none";
defparam ram_block3a41.port_b_data_width = 1;
defparam ram_block3a41.port_b_first_address = 0;
defparam ram_block3a41.port_b_first_bit_number = 9;
defparam ram_block3a41.port_b_last_address = 8191;
defparam ram_block3a41.port_b_logical_ram_depth = 16384;
defparam ram_block3a41.port_b_logical_ram_width = 32;
defparam ram_block3a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_read_enable_clock = "clock1";
defparam ram_block3a41.port_b_write_enable_clock = "clock1";
defparam ram_block3a41.ram_block_type = "M9K";
defparam ram_block3a41.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y36_N0
cycloneive_ram_block ram_block3a9(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a9_PORTADATAOUT_bus),
	.portbdataout(ram_block3a9_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a9.clk0_core_clock_enable = "ena0";
defparam ram_block3a9.clk1_core_clock_enable = "ena1";
defparam ram_block3a9.data_interleave_offset_in_bits = 1;
defparam ram_block3a9.data_interleave_width_in_bits = 1;
defparam ram_block3a9.init_file = "meminit.hex";
defparam ram_block3a9.init_file_layout = "port_a";
defparam ram_block3a9.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a9.operation_mode = "bidir_dual_port";
defparam ram_block3a9.port_a_address_clear = "none";
defparam ram_block3a9.port_a_address_width = 13;
defparam ram_block3a9.port_a_byte_enable_clock = "none";
defparam ram_block3a9.port_a_data_out_clear = "none";
defparam ram_block3a9.port_a_data_out_clock = "none";
defparam ram_block3a9.port_a_data_width = 1;
defparam ram_block3a9.port_a_first_address = 0;
defparam ram_block3a9.port_a_first_bit_number = 9;
defparam ram_block3a9.port_a_last_address = 8191;
defparam ram_block3a9.port_a_logical_ram_depth = 16384;
defparam ram_block3a9.port_a_logical_ram_width = 32;
defparam ram_block3a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_address_clear = "none";
defparam ram_block3a9.port_b_address_clock = "clock1";
defparam ram_block3a9.port_b_address_width = 13;
defparam ram_block3a9.port_b_data_in_clock = "clock1";
defparam ram_block3a9.port_b_data_out_clear = "none";
defparam ram_block3a9.port_b_data_out_clock = "none";
defparam ram_block3a9.port_b_data_width = 1;
defparam ram_block3a9.port_b_first_address = 0;
defparam ram_block3a9.port_b_first_bit_number = 9;
defparam ram_block3a9.port_b_last_address = 8191;
defparam ram_block3a9.port_b_logical_ram_depth = 16384;
defparam ram_block3a9.port_b_logical_ram_width = 32;
defparam ram_block3a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_read_enable_clock = "clock1";
defparam ram_block3a9.port_b_write_enable_clock = "clock1";
defparam ram_block3a9.ram_block_type = "M9K";
defparam ram_block3a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220220080F;
// synopsys translate_on

// Location: M9K_X64_Y42_N0
cycloneive_ram_block ram_block3a42(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a42_PORTADATAOUT_bus),
	.portbdataout(ram_block3a42_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a42.clk0_core_clock_enable = "ena0";
defparam ram_block3a42.clk1_core_clock_enable = "ena1";
defparam ram_block3a42.data_interleave_offset_in_bits = 1;
defparam ram_block3a42.data_interleave_width_in_bits = 1;
defparam ram_block3a42.init_file = "meminit.hex";
defparam ram_block3a42.init_file_layout = "port_a";
defparam ram_block3a42.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a42.operation_mode = "bidir_dual_port";
defparam ram_block3a42.port_a_address_clear = "none";
defparam ram_block3a42.port_a_address_width = 13;
defparam ram_block3a42.port_a_byte_enable_clock = "none";
defparam ram_block3a42.port_a_data_out_clear = "none";
defparam ram_block3a42.port_a_data_out_clock = "none";
defparam ram_block3a42.port_a_data_width = 1;
defparam ram_block3a42.port_a_first_address = 0;
defparam ram_block3a42.port_a_first_bit_number = 10;
defparam ram_block3a42.port_a_last_address = 8191;
defparam ram_block3a42.port_a_logical_ram_depth = 16384;
defparam ram_block3a42.port_a_logical_ram_width = 32;
defparam ram_block3a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_address_clear = "none";
defparam ram_block3a42.port_b_address_clock = "clock1";
defparam ram_block3a42.port_b_address_width = 13;
defparam ram_block3a42.port_b_data_in_clock = "clock1";
defparam ram_block3a42.port_b_data_out_clear = "none";
defparam ram_block3a42.port_b_data_out_clock = "none";
defparam ram_block3a42.port_b_data_width = 1;
defparam ram_block3a42.port_b_first_address = 0;
defparam ram_block3a42.port_b_first_bit_number = 10;
defparam ram_block3a42.port_b_last_address = 8191;
defparam ram_block3a42.port_b_logical_ram_depth = 16384;
defparam ram_block3a42.port_b_logical_ram_width = 32;
defparam ram_block3a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_read_enable_clock = "clock1";
defparam ram_block3a42.port_b_write_enable_clock = "clock1";
defparam ram_block3a42.ram_block_type = "M9K";
defparam ram_block3a42.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y43_N0
cycloneive_ram_block ram_block3a10(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a10_PORTADATAOUT_bus),
	.portbdataout(ram_block3a10_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a10.clk0_core_clock_enable = "ena0";
defparam ram_block3a10.clk1_core_clock_enable = "ena1";
defparam ram_block3a10.data_interleave_offset_in_bits = 1;
defparam ram_block3a10.data_interleave_width_in_bits = 1;
defparam ram_block3a10.init_file = "meminit.hex";
defparam ram_block3a10.init_file_layout = "port_a";
defparam ram_block3a10.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a10.operation_mode = "bidir_dual_port";
defparam ram_block3a10.port_a_address_clear = "none";
defparam ram_block3a10.port_a_address_width = 13;
defparam ram_block3a10.port_a_byte_enable_clock = "none";
defparam ram_block3a10.port_a_data_out_clear = "none";
defparam ram_block3a10.port_a_data_out_clock = "none";
defparam ram_block3a10.port_a_data_width = 1;
defparam ram_block3a10.port_a_first_address = 0;
defparam ram_block3a10.port_a_first_bit_number = 10;
defparam ram_block3a10.port_a_last_address = 8191;
defparam ram_block3a10.port_a_logical_ram_depth = 16384;
defparam ram_block3a10.port_a_logical_ram_width = 32;
defparam ram_block3a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_address_clear = "none";
defparam ram_block3a10.port_b_address_clock = "clock1";
defparam ram_block3a10.port_b_address_width = 13;
defparam ram_block3a10.port_b_data_in_clock = "clock1";
defparam ram_block3a10.port_b_data_out_clear = "none";
defparam ram_block3a10.port_b_data_out_clock = "none";
defparam ram_block3a10.port_b_data_width = 1;
defparam ram_block3a10.port_b_first_address = 0;
defparam ram_block3a10.port_b_first_bit_number = 10;
defparam ram_block3a10.port_b_last_address = 8191;
defparam ram_block3a10.port_b_logical_ram_depth = 16384;
defparam ram_block3a10.port_b_logical_ram_width = 32;
defparam ram_block3a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_read_enable_clock = "clock1";
defparam ram_block3a10.port_b_write_enable_clock = "clock1";
defparam ram_block3a10.ram_block_type = "M9K";
defparam ram_block3a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002202300003;
// synopsys translate_on

// Location: M9K_X78_Y41_N0
cycloneive_ram_block ram_block3a43(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a43_PORTADATAOUT_bus),
	.portbdataout(ram_block3a43_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a43.clk0_core_clock_enable = "ena0";
defparam ram_block3a43.clk1_core_clock_enable = "ena1";
defparam ram_block3a43.data_interleave_offset_in_bits = 1;
defparam ram_block3a43.data_interleave_width_in_bits = 1;
defparam ram_block3a43.init_file = "meminit.hex";
defparam ram_block3a43.init_file_layout = "port_a";
defparam ram_block3a43.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a43.operation_mode = "bidir_dual_port";
defparam ram_block3a43.port_a_address_clear = "none";
defparam ram_block3a43.port_a_address_width = 13;
defparam ram_block3a43.port_a_byte_enable_clock = "none";
defparam ram_block3a43.port_a_data_out_clear = "none";
defparam ram_block3a43.port_a_data_out_clock = "none";
defparam ram_block3a43.port_a_data_width = 1;
defparam ram_block3a43.port_a_first_address = 0;
defparam ram_block3a43.port_a_first_bit_number = 11;
defparam ram_block3a43.port_a_last_address = 8191;
defparam ram_block3a43.port_a_logical_ram_depth = 16384;
defparam ram_block3a43.port_a_logical_ram_width = 32;
defparam ram_block3a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_address_clear = "none";
defparam ram_block3a43.port_b_address_clock = "clock1";
defparam ram_block3a43.port_b_address_width = 13;
defparam ram_block3a43.port_b_data_in_clock = "clock1";
defparam ram_block3a43.port_b_data_out_clear = "none";
defparam ram_block3a43.port_b_data_out_clock = "none";
defparam ram_block3a43.port_b_data_width = 1;
defparam ram_block3a43.port_b_first_address = 0;
defparam ram_block3a43.port_b_first_bit_number = 11;
defparam ram_block3a43.port_b_last_address = 8191;
defparam ram_block3a43.port_b_logical_ram_depth = 16384;
defparam ram_block3a43.port_b_logical_ram_width = 32;
defparam ram_block3a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_read_enable_clock = "clock1";
defparam ram_block3a43.port_b_write_enable_clock = "clock1";
defparam ram_block3a43.ram_block_type = "M9K";
defparam ram_block3a43.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y45_N0
cycloneive_ram_block ram_block3a11(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a11_PORTADATAOUT_bus),
	.portbdataout(ram_block3a11_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a11.clk0_core_clock_enable = "ena0";
defparam ram_block3a11.clk1_core_clock_enable = "ena1";
defparam ram_block3a11.data_interleave_offset_in_bits = 1;
defparam ram_block3a11.data_interleave_width_in_bits = 1;
defparam ram_block3a11.init_file = "meminit.hex";
defparam ram_block3a11.init_file_layout = "port_a";
defparam ram_block3a11.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a11.operation_mode = "bidir_dual_port";
defparam ram_block3a11.port_a_address_clear = "none";
defparam ram_block3a11.port_a_address_width = 13;
defparam ram_block3a11.port_a_byte_enable_clock = "none";
defparam ram_block3a11.port_a_data_out_clear = "none";
defparam ram_block3a11.port_a_data_out_clock = "none";
defparam ram_block3a11.port_a_data_width = 1;
defparam ram_block3a11.port_a_first_address = 0;
defparam ram_block3a11.port_a_first_bit_number = 11;
defparam ram_block3a11.port_a_last_address = 8191;
defparam ram_block3a11.port_a_logical_ram_depth = 16384;
defparam ram_block3a11.port_a_logical_ram_width = 32;
defparam ram_block3a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_address_clear = "none";
defparam ram_block3a11.port_b_address_clock = "clock1";
defparam ram_block3a11.port_b_address_width = 13;
defparam ram_block3a11.port_b_data_in_clock = "clock1";
defparam ram_block3a11.port_b_data_out_clear = "none";
defparam ram_block3a11.port_b_data_out_clock = "none";
defparam ram_block3a11.port_b_data_width = 1;
defparam ram_block3a11.port_b_first_address = 0;
defparam ram_block3a11.port_b_first_bit_number = 11;
defparam ram_block3a11.port_b_last_address = 8191;
defparam ram_block3a11.port_b_logical_ram_depth = 16384;
defparam ram_block3a11.port_b_logical_ram_width = 32;
defparam ram_block3a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_read_enable_clock = "clock1";
defparam ram_block3a11.port_b_write_enable_clock = "clock1";
defparam ram_block3a11.ram_block_type = "M9K";
defparam ram_block3a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210800265A2A2233;
// synopsys translate_on

// Location: M9K_X51_Y44_N0
cycloneive_ram_block ram_block3a44(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a44_PORTADATAOUT_bus),
	.portbdataout(ram_block3a44_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a44.clk0_core_clock_enable = "ena0";
defparam ram_block3a44.clk1_core_clock_enable = "ena1";
defparam ram_block3a44.data_interleave_offset_in_bits = 1;
defparam ram_block3a44.data_interleave_width_in_bits = 1;
defparam ram_block3a44.init_file = "meminit.hex";
defparam ram_block3a44.init_file_layout = "port_a";
defparam ram_block3a44.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a44.operation_mode = "bidir_dual_port";
defparam ram_block3a44.port_a_address_clear = "none";
defparam ram_block3a44.port_a_address_width = 13;
defparam ram_block3a44.port_a_byte_enable_clock = "none";
defparam ram_block3a44.port_a_data_out_clear = "none";
defparam ram_block3a44.port_a_data_out_clock = "none";
defparam ram_block3a44.port_a_data_width = 1;
defparam ram_block3a44.port_a_first_address = 0;
defparam ram_block3a44.port_a_first_bit_number = 12;
defparam ram_block3a44.port_a_last_address = 8191;
defparam ram_block3a44.port_a_logical_ram_depth = 16384;
defparam ram_block3a44.port_a_logical_ram_width = 32;
defparam ram_block3a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_address_clear = "none";
defparam ram_block3a44.port_b_address_clock = "clock1";
defparam ram_block3a44.port_b_address_width = 13;
defparam ram_block3a44.port_b_data_in_clock = "clock1";
defparam ram_block3a44.port_b_data_out_clear = "none";
defparam ram_block3a44.port_b_data_out_clock = "none";
defparam ram_block3a44.port_b_data_width = 1;
defparam ram_block3a44.port_b_first_address = 0;
defparam ram_block3a44.port_b_first_bit_number = 12;
defparam ram_block3a44.port_b_last_address = 8191;
defparam ram_block3a44.port_b_logical_ram_depth = 16384;
defparam ram_block3a44.port_b_logical_ram_width = 32;
defparam ram_block3a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_read_enable_clock = "clock1";
defparam ram_block3a44.port_b_write_enable_clock = "clock1";
defparam ram_block3a44.ram_block_type = "M9K";
defparam ram_block3a44.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y47_N0
cycloneive_ram_block ram_block3a12(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a12_PORTADATAOUT_bus),
	.portbdataout(ram_block3a12_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a12.clk0_core_clock_enable = "ena0";
defparam ram_block3a12.clk1_core_clock_enable = "ena1";
defparam ram_block3a12.data_interleave_offset_in_bits = 1;
defparam ram_block3a12.data_interleave_width_in_bits = 1;
defparam ram_block3a12.init_file = "meminit.hex";
defparam ram_block3a12.init_file_layout = "port_a";
defparam ram_block3a12.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a12.operation_mode = "bidir_dual_port";
defparam ram_block3a12.port_a_address_clear = "none";
defparam ram_block3a12.port_a_address_width = 13;
defparam ram_block3a12.port_a_byte_enable_clock = "none";
defparam ram_block3a12.port_a_data_out_clear = "none";
defparam ram_block3a12.port_a_data_out_clock = "none";
defparam ram_block3a12.port_a_data_width = 1;
defparam ram_block3a12.port_a_first_address = 0;
defparam ram_block3a12.port_a_first_bit_number = 12;
defparam ram_block3a12.port_a_last_address = 8191;
defparam ram_block3a12.port_a_logical_ram_depth = 16384;
defparam ram_block3a12.port_a_logical_ram_width = 32;
defparam ram_block3a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_address_clear = "none";
defparam ram_block3a12.port_b_address_clock = "clock1";
defparam ram_block3a12.port_b_address_width = 13;
defparam ram_block3a12.port_b_data_in_clock = "clock1";
defparam ram_block3a12.port_b_data_out_clear = "none";
defparam ram_block3a12.port_b_data_out_clock = "none";
defparam ram_block3a12.port_b_data_width = 1;
defparam ram_block3a12.port_b_first_address = 0;
defparam ram_block3a12.port_b_first_bit_number = 12;
defparam ram_block3a12.port_b_last_address = 8191;
defparam ram_block3a12.port_b_logical_ram_depth = 16384;
defparam ram_block3a12.port_b_logical_ram_width = 32;
defparam ram_block3a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_read_enable_clock = "clock1";
defparam ram_block3a12.port_b_write_enable_clock = "clock1";
defparam ram_block3a12.ram_block_type = "M9K";
defparam ram_block3a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022C2043;
// synopsys translate_on

// Location: M9K_X64_Y29_N0
cycloneive_ram_block ram_block3a45(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a45_PORTADATAOUT_bus),
	.portbdataout(ram_block3a45_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a45.clk0_core_clock_enable = "ena0";
defparam ram_block3a45.clk1_core_clock_enable = "ena1";
defparam ram_block3a45.data_interleave_offset_in_bits = 1;
defparam ram_block3a45.data_interleave_width_in_bits = 1;
defparam ram_block3a45.init_file = "meminit.hex";
defparam ram_block3a45.init_file_layout = "port_a";
defparam ram_block3a45.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a45.operation_mode = "bidir_dual_port";
defparam ram_block3a45.port_a_address_clear = "none";
defparam ram_block3a45.port_a_address_width = 13;
defparam ram_block3a45.port_a_byte_enable_clock = "none";
defparam ram_block3a45.port_a_data_out_clear = "none";
defparam ram_block3a45.port_a_data_out_clock = "none";
defparam ram_block3a45.port_a_data_width = 1;
defparam ram_block3a45.port_a_first_address = 0;
defparam ram_block3a45.port_a_first_bit_number = 13;
defparam ram_block3a45.port_a_last_address = 8191;
defparam ram_block3a45.port_a_logical_ram_depth = 16384;
defparam ram_block3a45.port_a_logical_ram_width = 32;
defparam ram_block3a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_address_clear = "none";
defparam ram_block3a45.port_b_address_clock = "clock1";
defparam ram_block3a45.port_b_address_width = 13;
defparam ram_block3a45.port_b_data_in_clock = "clock1";
defparam ram_block3a45.port_b_data_out_clear = "none";
defparam ram_block3a45.port_b_data_out_clock = "none";
defparam ram_block3a45.port_b_data_width = 1;
defparam ram_block3a45.port_b_first_address = 0;
defparam ram_block3a45.port_b_first_bit_number = 13;
defparam ram_block3a45.port_b_last_address = 8191;
defparam ram_block3a45.port_b_logical_ram_depth = 16384;
defparam ram_block3a45.port_b_logical_ram_width = 32;
defparam ram_block3a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_read_enable_clock = "clock1";
defparam ram_block3a45.port_b_write_enable_clock = "clock1";
defparam ram_block3a45.ram_block_type = "M9K";
defparam ram_block3a45.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y29_N0
cycloneive_ram_block ram_block3a13(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a13_PORTADATAOUT_bus),
	.portbdataout(ram_block3a13_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a13.clk0_core_clock_enable = "ena0";
defparam ram_block3a13.clk1_core_clock_enable = "ena1";
defparam ram_block3a13.data_interleave_offset_in_bits = 1;
defparam ram_block3a13.data_interleave_width_in_bits = 1;
defparam ram_block3a13.init_file = "meminit.hex";
defparam ram_block3a13.init_file_layout = "port_a";
defparam ram_block3a13.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a13.operation_mode = "bidir_dual_port";
defparam ram_block3a13.port_a_address_clear = "none";
defparam ram_block3a13.port_a_address_width = 13;
defparam ram_block3a13.port_a_byte_enable_clock = "none";
defparam ram_block3a13.port_a_data_out_clear = "none";
defparam ram_block3a13.port_a_data_out_clock = "none";
defparam ram_block3a13.port_a_data_width = 1;
defparam ram_block3a13.port_a_first_address = 0;
defparam ram_block3a13.port_a_first_bit_number = 13;
defparam ram_block3a13.port_a_last_address = 8191;
defparam ram_block3a13.port_a_logical_ram_depth = 16384;
defparam ram_block3a13.port_a_logical_ram_width = 32;
defparam ram_block3a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_address_clear = "none";
defparam ram_block3a13.port_b_address_clock = "clock1";
defparam ram_block3a13.port_b_address_width = 13;
defparam ram_block3a13.port_b_data_in_clock = "clock1";
defparam ram_block3a13.port_b_data_out_clear = "none";
defparam ram_block3a13.port_b_data_out_clock = "none";
defparam ram_block3a13.port_b_data_width = 1;
defparam ram_block3a13.port_b_first_address = 0;
defparam ram_block3a13.port_b_first_bit_number = 13;
defparam ram_block3a13.port_b_last_address = 8191;
defparam ram_block3a13.port_b_logical_ram_depth = 16384;
defparam ram_block3a13.port_b_logical_ram_width = 32;
defparam ram_block3a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_read_enable_clock = "clock1";
defparam ram_block3a13.port_b_write_enable_clock = "clock1";
defparam ram_block3a13.ram_block_type = "M9K";
defparam ram_block3a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022F5213;
// synopsys translate_on

// Location: M9K_X64_Y28_N0
cycloneive_ram_block ram_block3a46(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a46_PORTADATAOUT_bus),
	.portbdataout(ram_block3a46_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a46.clk0_core_clock_enable = "ena0";
defparam ram_block3a46.clk1_core_clock_enable = "ena1";
defparam ram_block3a46.data_interleave_offset_in_bits = 1;
defparam ram_block3a46.data_interleave_width_in_bits = 1;
defparam ram_block3a46.init_file = "meminit.hex";
defparam ram_block3a46.init_file_layout = "port_a";
defparam ram_block3a46.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a46.operation_mode = "bidir_dual_port";
defparam ram_block3a46.port_a_address_clear = "none";
defparam ram_block3a46.port_a_address_width = 13;
defparam ram_block3a46.port_a_byte_enable_clock = "none";
defparam ram_block3a46.port_a_data_out_clear = "none";
defparam ram_block3a46.port_a_data_out_clock = "none";
defparam ram_block3a46.port_a_data_width = 1;
defparam ram_block3a46.port_a_first_address = 0;
defparam ram_block3a46.port_a_first_bit_number = 14;
defparam ram_block3a46.port_a_last_address = 8191;
defparam ram_block3a46.port_a_logical_ram_depth = 16384;
defparam ram_block3a46.port_a_logical_ram_width = 32;
defparam ram_block3a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_address_clear = "none";
defparam ram_block3a46.port_b_address_clock = "clock1";
defparam ram_block3a46.port_b_address_width = 13;
defparam ram_block3a46.port_b_data_in_clock = "clock1";
defparam ram_block3a46.port_b_data_out_clear = "none";
defparam ram_block3a46.port_b_data_out_clock = "none";
defparam ram_block3a46.port_b_data_width = 1;
defparam ram_block3a46.port_b_first_address = 0;
defparam ram_block3a46.port_b_first_bit_number = 14;
defparam ram_block3a46.port_b_last_address = 8191;
defparam ram_block3a46.port_b_logical_ram_depth = 16384;
defparam ram_block3a46.port_b_logical_ram_width = 32;
defparam ram_block3a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_read_enable_clock = "clock1";
defparam ram_block3a46.port_b_write_enable_clock = "clock1";
defparam ram_block3a46.ram_block_type = "M9K";
defparam ram_block3a46.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y33_N0
cycloneive_ram_block ram_block3a14(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a14_PORTADATAOUT_bus),
	.portbdataout(ram_block3a14_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a14.clk0_core_clock_enable = "ena0";
defparam ram_block3a14.clk1_core_clock_enable = "ena1";
defparam ram_block3a14.data_interleave_offset_in_bits = 1;
defparam ram_block3a14.data_interleave_width_in_bits = 1;
defparam ram_block3a14.init_file = "meminit.hex";
defparam ram_block3a14.init_file_layout = "port_a";
defparam ram_block3a14.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a14.operation_mode = "bidir_dual_port";
defparam ram_block3a14.port_a_address_clear = "none";
defparam ram_block3a14.port_a_address_width = 13;
defparam ram_block3a14.port_a_byte_enable_clock = "none";
defparam ram_block3a14.port_a_data_out_clear = "none";
defparam ram_block3a14.port_a_data_out_clock = "none";
defparam ram_block3a14.port_a_data_width = 1;
defparam ram_block3a14.port_a_first_address = 0;
defparam ram_block3a14.port_a_first_bit_number = 14;
defparam ram_block3a14.port_a_last_address = 8191;
defparam ram_block3a14.port_a_logical_ram_depth = 16384;
defparam ram_block3a14.port_a_logical_ram_width = 32;
defparam ram_block3a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_address_clear = "none";
defparam ram_block3a14.port_b_address_clock = "clock1";
defparam ram_block3a14.port_b_address_width = 13;
defparam ram_block3a14.port_b_data_in_clock = "clock1";
defparam ram_block3a14.port_b_data_out_clear = "none";
defparam ram_block3a14.port_b_data_out_clock = "none";
defparam ram_block3a14.port_b_data_width = 1;
defparam ram_block3a14.port_b_first_address = 0;
defparam ram_block3a14.port_b_first_bit_number = 14;
defparam ram_block3a14.port_b_last_address = 8191;
defparam ram_block3a14.port_b_logical_ram_depth = 16384;
defparam ram_block3a14.port_b_logical_ram_width = 32;
defparam ram_block3a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_read_enable_clock = "clock1";
defparam ram_block3a14.port_b_write_enable_clock = "clock1";
defparam ram_block3a14.ram_block_type = "M9K";
defparam ram_block3a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000224A200503;
// synopsys translate_on

// Location: M9K_X64_Y38_N0
cycloneive_ram_block ram_block3a47(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a47_PORTADATAOUT_bus),
	.portbdataout(ram_block3a47_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a47.clk0_core_clock_enable = "ena0";
defparam ram_block3a47.clk1_core_clock_enable = "ena1";
defparam ram_block3a47.data_interleave_offset_in_bits = 1;
defparam ram_block3a47.data_interleave_width_in_bits = 1;
defparam ram_block3a47.init_file = "meminit.hex";
defparam ram_block3a47.init_file_layout = "port_a";
defparam ram_block3a47.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a47.operation_mode = "bidir_dual_port";
defparam ram_block3a47.port_a_address_clear = "none";
defparam ram_block3a47.port_a_address_width = 13;
defparam ram_block3a47.port_a_byte_enable_clock = "none";
defparam ram_block3a47.port_a_data_out_clear = "none";
defparam ram_block3a47.port_a_data_out_clock = "none";
defparam ram_block3a47.port_a_data_width = 1;
defparam ram_block3a47.port_a_first_address = 0;
defparam ram_block3a47.port_a_first_bit_number = 15;
defparam ram_block3a47.port_a_last_address = 8191;
defparam ram_block3a47.port_a_logical_ram_depth = 16384;
defparam ram_block3a47.port_a_logical_ram_width = 32;
defparam ram_block3a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_address_clear = "none";
defparam ram_block3a47.port_b_address_clock = "clock1";
defparam ram_block3a47.port_b_address_width = 13;
defparam ram_block3a47.port_b_data_in_clock = "clock1";
defparam ram_block3a47.port_b_data_out_clear = "none";
defparam ram_block3a47.port_b_data_out_clock = "none";
defparam ram_block3a47.port_b_data_width = 1;
defparam ram_block3a47.port_b_first_address = 0;
defparam ram_block3a47.port_b_first_bit_number = 15;
defparam ram_block3a47.port_b_last_address = 8191;
defparam ram_block3a47.port_b_logical_ram_depth = 16384;
defparam ram_block3a47.port_b_logical_ram_width = 32;
defparam ram_block3a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_read_enable_clock = "clock1";
defparam ram_block3a47.port_b_write_enable_clock = "clock1";
defparam ram_block3a47.ram_block_type = "M9K";
defparam ram_block3a47.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y37_N0
cycloneive_ram_block ram_block3a15(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a15_PORTADATAOUT_bus),
	.portbdataout(ram_block3a15_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a15.clk0_core_clock_enable = "ena0";
defparam ram_block3a15.clk1_core_clock_enable = "ena1";
defparam ram_block3a15.data_interleave_offset_in_bits = 1;
defparam ram_block3a15.data_interleave_width_in_bits = 1;
defparam ram_block3a15.init_file = "meminit.hex";
defparam ram_block3a15.init_file_layout = "port_a";
defparam ram_block3a15.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a15.operation_mode = "bidir_dual_port";
defparam ram_block3a15.port_a_address_clear = "none";
defparam ram_block3a15.port_a_address_width = 13;
defparam ram_block3a15.port_a_byte_enable_clock = "none";
defparam ram_block3a15.port_a_data_out_clear = "none";
defparam ram_block3a15.port_a_data_out_clock = "none";
defparam ram_block3a15.port_a_data_width = 1;
defparam ram_block3a15.port_a_first_address = 0;
defparam ram_block3a15.port_a_first_bit_number = 15;
defparam ram_block3a15.port_a_last_address = 8191;
defparam ram_block3a15.port_a_logical_ram_depth = 16384;
defparam ram_block3a15.port_a_logical_ram_width = 32;
defparam ram_block3a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_address_clear = "none";
defparam ram_block3a15.port_b_address_clock = "clock1";
defparam ram_block3a15.port_b_address_width = 13;
defparam ram_block3a15.port_b_data_in_clock = "clock1";
defparam ram_block3a15.port_b_data_out_clear = "none";
defparam ram_block3a15.port_b_data_out_clock = "none";
defparam ram_block3a15.port_b_data_width = 1;
defparam ram_block3a15.port_b_first_address = 0;
defparam ram_block3a15.port_b_first_bit_number = 15;
defparam ram_block3a15.port_b_last_address = 8191;
defparam ram_block3a15.port_b_logical_ram_depth = 16384;
defparam ram_block3a15.port_b_logical_ram_width = 32;
defparam ram_block3a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_read_enable_clock = "clock1";
defparam ram_block3a15.port_b_write_enable_clock = "clock1";
defparam ram_block3a15.ram_block_type = "M9K";
defparam ram_block3a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002242206063;
// synopsys translate_on

// Location: M9K_X51_Y39_N0
cycloneive_ram_block ram_block3a48(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a48_PORTADATAOUT_bus),
	.portbdataout(ram_block3a48_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a48.clk0_core_clock_enable = "ena0";
defparam ram_block3a48.clk1_core_clock_enable = "ena1";
defparam ram_block3a48.data_interleave_offset_in_bits = 1;
defparam ram_block3a48.data_interleave_width_in_bits = 1;
defparam ram_block3a48.init_file = "meminit.hex";
defparam ram_block3a48.init_file_layout = "port_a";
defparam ram_block3a48.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a48.operation_mode = "bidir_dual_port";
defparam ram_block3a48.port_a_address_clear = "none";
defparam ram_block3a48.port_a_address_width = 13;
defparam ram_block3a48.port_a_byte_enable_clock = "none";
defparam ram_block3a48.port_a_data_out_clear = "none";
defparam ram_block3a48.port_a_data_out_clock = "none";
defparam ram_block3a48.port_a_data_width = 1;
defparam ram_block3a48.port_a_first_address = 0;
defparam ram_block3a48.port_a_first_bit_number = 16;
defparam ram_block3a48.port_a_last_address = 8191;
defparam ram_block3a48.port_a_logical_ram_depth = 16384;
defparam ram_block3a48.port_a_logical_ram_width = 32;
defparam ram_block3a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_address_clear = "none";
defparam ram_block3a48.port_b_address_clock = "clock1";
defparam ram_block3a48.port_b_address_width = 13;
defparam ram_block3a48.port_b_data_in_clock = "clock1";
defparam ram_block3a48.port_b_data_out_clear = "none";
defparam ram_block3a48.port_b_data_out_clock = "none";
defparam ram_block3a48.port_b_data_width = 1;
defparam ram_block3a48.port_b_first_address = 0;
defparam ram_block3a48.port_b_first_bit_number = 16;
defparam ram_block3a48.port_b_last_address = 8191;
defparam ram_block3a48.port_b_logical_ram_depth = 16384;
defparam ram_block3a48.port_b_logical_ram_width = 32;
defparam ram_block3a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_read_enable_clock = "clock1";
defparam ram_block3a48.port_b_write_enable_clock = "clock1";
defparam ram_block3a48.ram_block_type = "M9K";
defparam ram_block3a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y36_N0
cycloneive_ram_block ram_block3a16(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a16_PORTADATAOUT_bus),
	.portbdataout(ram_block3a16_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a16.clk0_core_clock_enable = "ena0";
defparam ram_block3a16.clk1_core_clock_enable = "ena1";
defparam ram_block3a16.data_interleave_offset_in_bits = 1;
defparam ram_block3a16.data_interleave_width_in_bits = 1;
defparam ram_block3a16.init_file = "meminit.hex";
defparam ram_block3a16.init_file_layout = "port_a";
defparam ram_block3a16.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a16.operation_mode = "bidir_dual_port";
defparam ram_block3a16.port_a_address_clear = "none";
defparam ram_block3a16.port_a_address_width = 13;
defparam ram_block3a16.port_a_byte_enable_clock = "none";
defparam ram_block3a16.port_a_data_out_clear = "none";
defparam ram_block3a16.port_a_data_out_clock = "none";
defparam ram_block3a16.port_a_data_width = 1;
defparam ram_block3a16.port_a_first_address = 0;
defparam ram_block3a16.port_a_first_bit_number = 16;
defparam ram_block3a16.port_a_last_address = 8191;
defparam ram_block3a16.port_a_logical_ram_depth = 16384;
defparam ram_block3a16.port_a_logical_ram_width = 32;
defparam ram_block3a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_address_clear = "none";
defparam ram_block3a16.port_b_address_clock = "clock1";
defparam ram_block3a16.port_b_address_width = 13;
defparam ram_block3a16.port_b_data_in_clock = "clock1";
defparam ram_block3a16.port_b_data_out_clear = "none";
defparam ram_block3a16.port_b_data_out_clock = "none";
defparam ram_block3a16.port_b_data_width = 1;
defparam ram_block3a16.port_b_first_address = 0;
defparam ram_block3a16.port_b_first_bit_number = 16;
defparam ram_block3a16.port_b_last_address = 8191;
defparam ram_block3a16.port_b_logical_ram_depth = 16384;
defparam ram_block3a16.port_b_logical_ram_width = 32;
defparam ram_block3a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_read_enable_clock = "clock1";
defparam ram_block3a16.port_b_write_enable_clock = "clock1";
defparam ram_block3a16.ram_block_type = "M9K";
defparam ram_block3a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000205A122003613254042;
// synopsys translate_on

// Location: M9K_X51_Y37_N0
cycloneive_ram_block ram_block3a49(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a49_PORTADATAOUT_bus),
	.portbdataout(ram_block3a49_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a49.clk0_core_clock_enable = "ena0";
defparam ram_block3a49.clk1_core_clock_enable = "ena1";
defparam ram_block3a49.data_interleave_offset_in_bits = 1;
defparam ram_block3a49.data_interleave_width_in_bits = 1;
defparam ram_block3a49.init_file = "meminit.hex";
defparam ram_block3a49.init_file_layout = "port_a";
defparam ram_block3a49.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a49.operation_mode = "bidir_dual_port";
defparam ram_block3a49.port_a_address_clear = "none";
defparam ram_block3a49.port_a_address_width = 13;
defparam ram_block3a49.port_a_byte_enable_clock = "none";
defparam ram_block3a49.port_a_data_out_clear = "none";
defparam ram_block3a49.port_a_data_out_clock = "none";
defparam ram_block3a49.port_a_data_width = 1;
defparam ram_block3a49.port_a_first_address = 0;
defparam ram_block3a49.port_a_first_bit_number = 17;
defparam ram_block3a49.port_a_last_address = 8191;
defparam ram_block3a49.port_a_logical_ram_depth = 16384;
defparam ram_block3a49.port_a_logical_ram_width = 32;
defparam ram_block3a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_address_clear = "none";
defparam ram_block3a49.port_b_address_clock = "clock1";
defparam ram_block3a49.port_b_address_width = 13;
defparam ram_block3a49.port_b_data_in_clock = "clock1";
defparam ram_block3a49.port_b_data_out_clear = "none";
defparam ram_block3a49.port_b_data_out_clock = "none";
defparam ram_block3a49.port_b_data_width = 1;
defparam ram_block3a49.port_b_first_address = 0;
defparam ram_block3a49.port_b_first_bit_number = 17;
defparam ram_block3a49.port_b_last_address = 8191;
defparam ram_block3a49.port_b_logical_ram_depth = 16384;
defparam ram_block3a49.port_b_logical_ram_width = 32;
defparam ram_block3a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_read_enable_clock = "clock1";
defparam ram_block3a49.port_b_write_enable_clock = "clock1";
defparam ram_block3a49.ram_block_type = "M9K";
defparam ram_block3a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y33_N0
cycloneive_ram_block ram_block3a17(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a17_PORTADATAOUT_bus),
	.portbdataout(ram_block3a17_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a17.clk0_core_clock_enable = "ena0";
defparam ram_block3a17.clk1_core_clock_enable = "ena1";
defparam ram_block3a17.data_interleave_offset_in_bits = 1;
defparam ram_block3a17.data_interleave_width_in_bits = 1;
defparam ram_block3a17.init_file = "meminit.hex";
defparam ram_block3a17.init_file_layout = "port_a";
defparam ram_block3a17.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a17.operation_mode = "bidir_dual_port";
defparam ram_block3a17.port_a_address_clear = "none";
defparam ram_block3a17.port_a_address_width = 13;
defparam ram_block3a17.port_a_byte_enable_clock = "none";
defparam ram_block3a17.port_a_data_out_clear = "none";
defparam ram_block3a17.port_a_data_out_clock = "none";
defparam ram_block3a17.port_a_data_width = 1;
defparam ram_block3a17.port_a_first_address = 0;
defparam ram_block3a17.port_a_first_bit_number = 17;
defparam ram_block3a17.port_a_last_address = 8191;
defparam ram_block3a17.port_a_logical_ram_depth = 16384;
defparam ram_block3a17.port_a_logical_ram_width = 32;
defparam ram_block3a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_address_clear = "none";
defparam ram_block3a17.port_b_address_clock = "clock1";
defparam ram_block3a17.port_b_address_width = 13;
defparam ram_block3a17.port_b_data_in_clock = "clock1";
defparam ram_block3a17.port_b_data_out_clear = "none";
defparam ram_block3a17.port_b_data_out_clock = "none";
defparam ram_block3a17.port_b_data_width = 1;
defparam ram_block3a17.port_b_first_address = 0;
defparam ram_block3a17.port_b_first_bit_number = 17;
defparam ram_block3a17.port_b_last_address = 8191;
defparam ram_block3a17.port_b_logical_ram_depth = 16384;
defparam ram_block3a17.port_b_logical_ram_width = 32;
defparam ram_block3a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_read_enable_clock = "clock1";
defparam ram_block3a17.port_b_write_enable_clock = "clock1";
defparam ram_block3a17.ram_block_type = "M9K";
defparam ram_block3a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006C0340C001602060001;
// synopsys translate_on

// Location: M9K_X37_Y37_N0
cycloneive_ram_block ram_block3a50(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a50_PORTADATAOUT_bus),
	.portbdataout(ram_block3a50_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a50.clk0_core_clock_enable = "ena0";
defparam ram_block3a50.clk1_core_clock_enable = "ena1";
defparam ram_block3a50.data_interleave_offset_in_bits = 1;
defparam ram_block3a50.data_interleave_width_in_bits = 1;
defparam ram_block3a50.init_file = "meminit.hex";
defparam ram_block3a50.init_file_layout = "port_a";
defparam ram_block3a50.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a50.operation_mode = "bidir_dual_port";
defparam ram_block3a50.port_a_address_clear = "none";
defparam ram_block3a50.port_a_address_width = 13;
defparam ram_block3a50.port_a_byte_enable_clock = "none";
defparam ram_block3a50.port_a_data_out_clear = "none";
defparam ram_block3a50.port_a_data_out_clock = "none";
defparam ram_block3a50.port_a_data_width = 1;
defparam ram_block3a50.port_a_first_address = 0;
defparam ram_block3a50.port_a_first_bit_number = 18;
defparam ram_block3a50.port_a_last_address = 8191;
defparam ram_block3a50.port_a_logical_ram_depth = 16384;
defparam ram_block3a50.port_a_logical_ram_width = 32;
defparam ram_block3a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_address_clear = "none";
defparam ram_block3a50.port_b_address_clock = "clock1";
defparam ram_block3a50.port_b_address_width = 13;
defparam ram_block3a50.port_b_data_in_clock = "clock1";
defparam ram_block3a50.port_b_data_out_clear = "none";
defparam ram_block3a50.port_b_data_out_clock = "none";
defparam ram_block3a50.port_b_data_width = 1;
defparam ram_block3a50.port_b_first_address = 0;
defparam ram_block3a50.port_b_first_bit_number = 18;
defparam ram_block3a50.port_b_last_address = 8191;
defparam ram_block3a50.port_b_logical_ram_depth = 16384;
defparam ram_block3a50.port_b_logical_ram_width = 32;
defparam ram_block3a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_read_enable_clock = "clock1";
defparam ram_block3a50.port_b_write_enable_clock = "clock1";
defparam ram_block3a50.ram_block_type = "M9K";
defparam ram_block3a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y37_N0
cycloneive_ram_block ram_block3a18(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a18_PORTADATAOUT_bus),
	.portbdataout(ram_block3a18_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a18.clk0_core_clock_enable = "ena0";
defparam ram_block3a18.clk1_core_clock_enable = "ena1";
defparam ram_block3a18.data_interleave_offset_in_bits = 1;
defparam ram_block3a18.data_interleave_width_in_bits = 1;
defparam ram_block3a18.init_file = "meminit.hex";
defparam ram_block3a18.init_file_layout = "port_a";
defparam ram_block3a18.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a18.operation_mode = "bidir_dual_port";
defparam ram_block3a18.port_a_address_clear = "none";
defparam ram_block3a18.port_a_address_width = 13;
defparam ram_block3a18.port_a_byte_enable_clock = "none";
defparam ram_block3a18.port_a_data_out_clear = "none";
defparam ram_block3a18.port_a_data_out_clock = "none";
defparam ram_block3a18.port_a_data_width = 1;
defparam ram_block3a18.port_a_first_address = 0;
defparam ram_block3a18.port_a_first_bit_number = 18;
defparam ram_block3a18.port_a_last_address = 8191;
defparam ram_block3a18.port_a_logical_ram_depth = 16384;
defparam ram_block3a18.port_a_logical_ram_width = 32;
defparam ram_block3a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_address_clear = "none";
defparam ram_block3a18.port_b_address_clock = "clock1";
defparam ram_block3a18.port_b_address_width = 13;
defparam ram_block3a18.port_b_data_in_clock = "clock1";
defparam ram_block3a18.port_b_data_out_clear = "none";
defparam ram_block3a18.port_b_data_out_clock = "none";
defparam ram_block3a18.port_b_data_width = 1;
defparam ram_block3a18.port_b_first_address = 0;
defparam ram_block3a18.port_b_first_bit_number = 18;
defparam ram_block3a18.port_b_last_address = 8191;
defparam ram_block3a18.port_b_logical_ram_depth = 16384;
defparam ram_block3a18.port_b_logical_ram_width = 32;
defparam ram_block3a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_read_enable_clock = "clock1";
defparam ram_block3a18.port_b_write_enable_clock = "clock1";
defparam ram_block3a18.ram_block_type = "M9K";
defparam ram_block3a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060C3180001703286867;
// synopsys translate_on

// Location: M9K_X64_Y32_N0
cycloneive_ram_block ram_block3a51(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a51_PORTADATAOUT_bus),
	.portbdataout(ram_block3a51_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a51.clk0_core_clock_enable = "ena0";
defparam ram_block3a51.clk1_core_clock_enable = "ena1";
defparam ram_block3a51.data_interleave_offset_in_bits = 1;
defparam ram_block3a51.data_interleave_width_in_bits = 1;
defparam ram_block3a51.init_file = "meminit.hex";
defparam ram_block3a51.init_file_layout = "port_a";
defparam ram_block3a51.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a51.operation_mode = "bidir_dual_port";
defparam ram_block3a51.port_a_address_clear = "none";
defparam ram_block3a51.port_a_address_width = 13;
defparam ram_block3a51.port_a_byte_enable_clock = "none";
defparam ram_block3a51.port_a_data_out_clear = "none";
defparam ram_block3a51.port_a_data_out_clock = "none";
defparam ram_block3a51.port_a_data_width = 1;
defparam ram_block3a51.port_a_first_address = 0;
defparam ram_block3a51.port_a_first_bit_number = 19;
defparam ram_block3a51.port_a_last_address = 8191;
defparam ram_block3a51.port_a_logical_ram_depth = 16384;
defparam ram_block3a51.port_a_logical_ram_width = 32;
defparam ram_block3a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_address_clear = "none";
defparam ram_block3a51.port_b_address_clock = "clock1";
defparam ram_block3a51.port_b_address_width = 13;
defparam ram_block3a51.port_b_data_in_clock = "clock1";
defparam ram_block3a51.port_b_data_out_clear = "none";
defparam ram_block3a51.port_b_data_out_clock = "none";
defparam ram_block3a51.port_b_data_width = 1;
defparam ram_block3a51.port_b_first_address = 0;
defparam ram_block3a51.port_b_first_bit_number = 19;
defparam ram_block3a51.port_b_last_address = 8191;
defparam ram_block3a51.port_b_logical_ram_depth = 16384;
defparam ram_block3a51.port_b_logical_ram_width = 32;
defparam ram_block3a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_read_enable_clock = "clock1";
defparam ram_block3a51.port_b_write_enable_clock = "clock1";
defparam ram_block3a51.ram_block_type = "M9K";
defparam ram_block3a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y33_N0
cycloneive_ram_block ram_block3a19(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a19_PORTADATAOUT_bus),
	.portbdataout(ram_block3a19_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a19.clk0_core_clock_enable = "ena0";
defparam ram_block3a19.clk1_core_clock_enable = "ena1";
defparam ram_block3a19.data_interleave_offset_in_bits = 1;
defparam ram_block3a19.data_interleave_width_in_bits = 1;
defparam ram_block3a19.init_file = "meminit.hex";
defparam ram_block3a19.init_file_layout = "port_a";
defparam ram_block3a19.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a19.operation_mode = "bidir_dual_port";
defparam ram_block3a19.port_a_address_clear = "none";
defparam ram_block3a19.port_a_address_width = 13;
defparam ram_block3a19.port_a_byte_enable_clock = "none";
defparam ram_block3a19.port_a_data_out_clear = "none";
defparam ram_block3a19.port_a_data_out_clock = "none";
defparam ram_block3a19.port_a_data_width = 1;
defparam ram_block3a19.port_a_first_address = 0;
defparam ram_block3a19.port_a_first_bit_number = 19;
defparam ram_block3a19.port_a_last_address = 8191;
defparam ram_block3a19.port_a_logical_ram_depth = 16384;
defparam ram_block3a19.port_a_logical_ram_width = 32;
defparam ram_block3a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_address_clear = "none";
defparam ram_block3a19.port_b_address_clock = "clock1";
defparam ram_block3a19.port_b_address_width = 13;
defparam ram_block3a19.port_b_data_in_clock = "clock1";
defparam ram_block3a19.port_b_data_out_clear = "none";
defparam ram_block3a19.port_b_data_out_clock = "none";
defparam ram_block3a19.port_b_data_width = 1;
defparam ram_block3a19.port_b_first_address = 0;
defparam ram_block3a19.port_b_first_bit_number = 19;
defparam ram_block3a19.port_b_last_address = 8191;
defparam ram_block3a19.port_b_logical_ram_depth = 16384;
defparam ram_block3a19.port_b_logical_ram_width = 32;
defparam ram_block3a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_read_enable_clock = "clock1";
defparam ram_block3a19.port_b_write_enable_clock = "clock1";
defparam ram_block3a19.ram_block_type = "M9K";
defparam ram_block3a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001C38C6E09B6D7701203;
// synopsys translate_on

// Location: M9K_X64_Y34_N0
cycloneive_ram_block ram_block3a52(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a52_PORTADATAOUT_bus),
	.portbdataout(ram_block3a52_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a52.clk0_core_clock_enable = "ena0";
defparam ram_block3a52.clk1_core_clock_enable = "ena1";
defparam ram_block3a52.data_interleave_offset_in_bits = 1;
defparam ram_block3a52.data_interleave_width_in_bits = 1;
defparam ram_block3a52.init_file = "meminit.hex";
defparam ram_block3a52.init_file_layout = "port_a";
defparam ram_block3a52.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a52.operation_mode = "bidir_dual_port";
defparam ram_block3a52.port_a_address_clear = "none";
defparam ram_block3a52.port_a_address_width = 13;
defparam ram_block3a52.port_a_byte_enable_clock = "none";
defparam ram_block3a52.port_a_data_out_clear = "none";
defparam ram_block3a52.port_a_data_out_clock = "none";
defparam ram_block3a52.port_a_data_width = 1;
defparam ram_block3a52.port_a_first_address = 0;
defparam ram_block3a52.port_a_first_bit_number = 20;
defparam ram_block3a52.port_a_last_address = 8191;
defparam ram_block3a52.port_a_logical_ram_depth = 16384;
defparam ram_block3a52.port_a_logical_ram_width = 32;
defparam ram_block3a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_address_clear = "none";
defparam ram_block3a52.port_b_address_clock = "clock1";
defparam ram_block3a52.port_b_address_width = 13;
defparam ram_block3a52.port_b_data_in_clock = "clock1";
defparam ram_block3a52.port_b_data_out_clear = "none";
defparam ram_block3a52.port_b_data_out_clock = "none";
defparam ram_block3a52.port_b_data_width = 1;
defparam ram_block3a52.port_b_first_address = 0;
defparam ram_block3a52.port_b_first_bit_number = 20;
defparam ram_block3a52.port_b_last_address = 8191;
defparam ram_block3a52.port_b_logical_ram_depth = 16384;
defparam ram_block3a52.port_b_logical_ram_width = 32;
defparam ram_block3a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_read_enable_clock = "clock1";
defparam ram_block3a52.port_b_write_enable_clock = "clock1";
defparam ram_block3a52.ram_block_type = "M9K";
defparam ram_block3a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y45_N0
cycloneive_ram_block ram_block3a20(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a20_PORTADATAOUT_bus),
	.portbdataout(ram_block3a20_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a20.clk0_core_clock_enable = "ena0";
defparam ram_block3a20.clk1_core_clock_enable = "ena1";
defparam ram_block3a20.data_interleave_offset_in_bits = 1;
defparam ram_block3a20.data_interleave_width_in_bits = 1;
defparam ram_block3a20.init_file = "meminit.hex";
defparam ram_block3a20.init_file_layout = "port_a";
defparam ram_block3a20.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a20.operation_mode = "bidir_dual_port";
defparam ram_block3a20.port_a_address_clear = "none";
defparam ram_block3a20.port_a_address_width = 13;
defparam ram_block3a20.port_a_byte_enable_clock = "none";
defparam ram_block3a20.port_a_data_out_clear = "none";
defparam ram_block3a20.port_a_data_out_clock = "none";
defparam ram_block3a20.port_a_data_width = 1;
defparam ram_block3a20.port_a_first_address = 0;
defparam ram_block3a20.port_a_first_bit_number = 20;
defparam ram_block3a20.port_a_last_address = 8191;
defparam ram_block3a20.port_a_logical_ram_depth = 16384;
defparam ram_block3a20.port_a_logical_ram_width = 32;
defparam ram_block3a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_address_clear = "none";
defparam ram_block3a20.port_b_address_clock = "clock1";
defparam ram_block3a20.port_b_address_width = 13;
defparam ram_block3a20.port_b_data_in_clock = "clock1";
defparam ram_block3a20.port_b_data_out_clear = "none";
defparam ram_block3a20.port_b_data_out_clock = "none";
defparam ram_block3a20.port_b_data_width = 1;
defparam ram_block3a20.port_b_first_address = 0;
defparam ram_block3a20.port_b_first_bit_number = 20;
defparam ram_block3a20.port_b_last_address = 8191;
defparam ram_block3a20.port_b_logical_ram_depth = 16384;
defparam ram_block3a20.port_b_logical_ram_width = 32;
defparam ram_block3a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_read_enable_clock = "clock1";
defparam ram_block3a20.port_b_write_enable_clock = "clock1";
defparam ram_block3a20.ram_block_type = "M9K";
defparam ram_block3a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A0832F000B;
// synopsys translate_on

// Location: M9K_X51_Y40_N0
cycloneive_ram_block ram_block3a53(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a53_PORTADATAOUT_bus),
	.portbdataout(ram_block3a53_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a53.clk0_core_clock_enable = "ena0";
defparam ram_block3a53.clk1_core_clock_enable = "ena1";
defparam ram_block3a53.data_interleave_offset_in_bits = 1;
defparam ram_block3a53.data_interleave_width_in_bits = 1;
defparam ram_block3a53.init_file = "meminit.hex";
defparam ram_block3a53.init_file_layout = "port_a";
defparam ram_block3a53.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a53.operation_mode = "bidir_dual_port";
defparam ram_block3a53.port_a_address_clear = "none";
defparam ram_block3a53.port_a_address_width = 13;
defparam ram_block3a53.port_a_byte_enable_clock = "none";
defparam ram_block3a53.port_a_data_out_clear = "none";
defparam ram_block3a53.port_a_data_out_clock = "none";
defparam ram_block3a53.port_a_data_width = 1;
defparam ram_block3a53.port_a_first_address = 0;
defparam ram_block3a53.port_a_first_bit_number = 21;
defparam ram_block3a53.port_a_last_address = 8191;
defparam ram_block3a53.port_a_logical_ram_depth = 16384;
defparam ram_block3a53.port_a_logical_ram_width = 32;
defparam ram_block3a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_address_clear = "none";
defparam ram_block3a53.port_b_address_clock = "clock1";
defparam ram_block3a53.port_b_address_width = 13;
defparam ram_block3a53.port_b_data_in_clock = "clock1";
defparam ram_block3a53.port_b_data_out_clear = "none";
defparam ram_block3a53.port_b_data_out_clock = "none";
defparam ram_block3a53.port_b_data_width = 1;
defparam ram_block3a53.port_b_first_address = 0;
defparam ram_block3a53.port_b_first_bit_number = 21;
defparam ram_block3a53.port_b_last_address = 8191;
defparam ram_block3a53.port_b_logical_ram_depth = 16384;
defparam ram_block3a53.port_b_logical_ram_width = 32;
defparam ram_block3a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_read_enable_clock = "clock1";
defparam ram_block3a53.port_b_write_enable_clock = "clock1";
defparam ram_block3a53.ram_block_type = "M9K";
defparam ram_block3a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y41_N0
cycloneive_ram_block ram_block3a21(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a21_PORTADATAOUT_bus),
	.portbdataout(ram_block3a21_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a21.clk0_core_clock_enable = "ena0";
defparam ram_block3a21.clk1_core_clock_enable = "ena1";
defparam ram_block3a21.data_interleave_offset_in_bits = 1;
defparam ram_block3a21.data_interleave_width_in_bits = 1;
defparam ram_block3a21.init_file = "meminit.hex";
defparam ram_block3a21.init_file_layout = "port_a";
defparam ram_block3a21.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a21.operation_mode = "bidir_dual_port";
defparam ram_block3a21.port_a_address_clear = "none";
defparam ram_block3a21.port_a_address_width = 13;
defparam ram_block3a21.port_a_byte_enable_clock = "none";
defparam ram_block3a21.port_a_data_out_clear = "none";
defparam ram_block3a21.port_a_data_out_clock = "none";
defparam ram_block3a21.port_a_data_width = 1;
defparam ram_block3a21.port_a_first_address = 0;
defparam ram_block3a21.port_a_first_bit_number = 21;
defparam ram_block3a21.port_a_last_address = 8191;
defparam ram_block3a21.port_a_logical_ram_depth = 16384;
defparam ram_block3a21.port_a_logical_ram_width = 32;
defparam ram_block3a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_address_clear = "none";
defparam ram_block3a21.port_b_address_clock = "clock1";
defparam ram_block3a21.port_b_address_width = 13;
defparam ram_block3a21.port_b_data_in_clock = "clock1";
defparam ram_block3a21.port_b_data_out_clear = "none";
defparam ram_block3a21.port_b_data_out_clock = "none";
defparam ram_block3a21.port_b_data_width = 1;
defparam ram_block3a21.port_b_first_address = 0;
defparam ram_block3a21.port_b_first_bit_number = 21;
defparam ram_block3a21.port_b_last_address = 8191;
defparam ram_block3a21.port_b_logical_ram_depth = 16384;
defparam ram_block3a21.port_b_logical_ram_width = 32;
defparam ram_block3a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_read_enable_clock = "clock1";
defparam ram_block3a21.port_b_write_enable_clock = "clock1";
defparam ram_block3a21.ram_block_type = "M9K";
defparam ram_block3a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002A142119BCBBAB600000;
// synopsys translate_on

// Location: M9K_X64_Y35_N0
cycloneive_ram_block ram_block3a54(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a54_PORTADATAOUT_bus),
	.portbdataout(ram_block3a54_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a54.clk0_core_clock_enable = "ena0";
defparam ram_block3a54.clk1_core_clock_enable = "ena1";
defparam ram_block3a54.data_interleave_offset_in_bits = 1;
defparam ram_block3a54.data_interleave_width_in_bits = 1;
defparam ram_block3a54.init_file = "meminit.hex";
defparam ram_block3a54.init_file_layout = "port_a";
defparam ram_block3a54.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a54.operation_mode = "bidir_dual_port";
defparam ram_block3a54.port_a_address_clear = "none";
defparam ram_block3a54.port_a_address_width = 13;
defparam ram_block3a54.port_a_byte_enable_clock = "none";
defparam ram_block3a54.port_a_data_out_clear = "none";
defparam ram_block3a54.port_a_data_out_clock = "none";
defparam ram_block3a54.port_a_data_width = 1;
defparam ram_block3a54.port_a_first_address = 0;
defparam ram_block3a54.port_a_first_bit_number = 22;
defparam ram_block3a54.port_a_last_address = 8191;
defparam ram_block3a54.port_a_logical_ram_depth = 16384;
defparam ram_block3a54.port_a_logical_ram_width = 32;
defparam ram_block3a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_address_clear = "none";
defparam ram_block3a54.port_b_address_clock = "clock1";
defparam ram_block3a54.port_b_address_width = 13;
defparam ram_block3a54.port_b_data_in_clock = "clock1";
defparam ram_block3a54.port_b_data_out_clear = "none";
defparam ram_block3a54.port_b_data_out_clock = "none";
defparam ram_block3a54.port_b_data_width = 1;
defparam ram_block3a54.port_b_first_address = 0;
defparam ram_block3a54.port_b_first_bit_number = 22;
defparam ram_block3a54.port_b_last_address = 8191;
defparam ram_block3a54.port_b_logical_ram_depth = 16384;
defparam ram_block3a54.port_b_logical_ram_width = 32;
defparam ram_block3a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_read_enable_clock = "clock1";
defparam ram_block3a54.port_b_write_enable_clock = "clock1";
defparam ram_block3a54.ram_block_type = "M9K";
defparam ram_block3a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y35_N0
cycloneive_ram_block ram_block3a22(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a22_PORTADATAOUT_bus),
	.portbdataout(ram_block3a22_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a22.clk0_core_clock_enable = "ena0";
defparam ram_block3a22.clk1_core_clock_enable = "ena1";
defparam ram_block3a22.data_interleave_offset_in_bits = 1;
defparam ram_block3a22.data_interleave_width_in_bits = 1;
defparam ram_block3a22.init_file = "meminit.hex";
defparam ram_block3a22.init_file_layout = "port_a";
defparam ram_block3a22.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a22.operation_mode = "bidir_dual_port";
defparam ram_block3a22.port_a_address_clear = "none";
defparam ram_block3a22.port_a_address_width = 13;
defparam ram_block3a22.port_a_byte_enable_clock = "none";
defparam ram_block3a22.port_a_data_out_clear = "none";
defparam ram_block3a22.port_a_data_out_clock = "none";
defparam ram_block3a22.port_a_data_width = 1;
defparam ram_block3a22.port_a_first_address = 0;
defparam ram_block3a22.port_a_first_bit_number = 22;
defparam ram_block3a22.port_a_last_address = 8191;
defparam ram_block3a22.port_a_logical_ram_depth = 16384;
defparam ram_block3a22.port_a_logical_ram_width = 32;
defparam ram_block3a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_address_clear = "none";
defparam ram_block3a22.port_b_address_clock = "clock1";
defparam ram_block3a22.port_b_address_width = 13;
defparam ram_block3a22.port_b_data_in_clock = "clock1";
defparam ram_block3a22.port_b_data_out_clear = "none";
defparam ram_block3a22.port_b_data_out_clock = "none";
defparam ram_block3a22.port_b_data_width = 1;
defparam ram_block3a22.port_b_first_address = 0;
defparam ram_block3a22.port_b_first_bit_number = 22;
defparam ram_block3a22.port_b_last_address = 8191;
defparam ram_block3a22.port_b_logical_ram_depth = 16384;
defparam ram_block3a22.port_b_logical_ram_width = 32;
defparam ram_block3a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_read_enable_clock = "clock1";
defparam ram_block3a22.port_b_write_enable_clock = "clock1";
defparam ram_block3a22.ram_block_type = "M9K";
defparam ram_block3a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E403004A40002000000;
// synopsys translate_on

// Location: M9K_X51_Y34_N0
cycloneive_ram_block ram_block3a55(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a55_PORTADATAOUT_bus),
	.portbdataout(ram_block3a55_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a55.clk0_core_clock_enable = "ena0";
defparam ram_block3a55.clk1_core_clock_enable = "ena1";
defparam ram_block3a55.data_interleave_offset_in_bits = 1;
defparam ram_block3a55.data_interleave_width_in_bits = 1;
defparam ram_block3a55.init_file = "meminit.hex";
defparam ram_block3a55.init_file_layout = "port_a";
defparam ram_block3a55.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a55.operation_mode = "bidir_dual_port";
defparam ram_block3a55.port_a_address_clear = "none";
defparam ram_block3a55.port_a_address_width = 13;
defparam ram_block3a55.port_a_byte_enable_clock = "none";
defparam ram_block3a55.port_a_data_out_clear = "none";
defparam ram_block3a55.port_a_data_out_clock = "none";
defparam ram_block3a55.port_a_data_width = 1;
defparam ram_block3a55.port_a_first_address = 0;
defparam ram_block3a55.port_a_first_bit_number = 23;
defparam ram_block3a55.port_a_last_address = 8191;
defparam ram_block3a55.port_a_logical_ram_depth = 16384;
defparam ram_block3a55.port_a_logical_ram_width = 32;
defparam ram_block3a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_address_clear = "none";
defparam ram_block3a55.port_b_address_clock = "clock1";
defparam ram_block3a55.port_b_address_width = 13;
defparam ram_block3a55.port_b_data_in_clock = "clock1";
defparam ram_block3a55.port_b_data_out_clear = "none";
defparam ram_block3a55.port_b_data_out_clock = "none";
defparam ram_block3a55.port_b_data_width = 1;
defparam ram_block3a55.port_b_first_address = 0;
defparam ram_block3a55.port_b_first_bit_number = 23;
defparam ram_block3a55.port_b_last_address = 8191;
defparam ram_block3a55.port_b_logical_ram_depth = 16384;
defparam ram_block3a55.port_b_logical_ram_width = 32;
defparam ram_block3a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_read_enable_clock = "clock1";
defparam ram_block3a55.port_b_write_enable_clock = "clock1";
defparam ram_block3a55.ram_block_type = "M9K";
defparam ram_block3a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y31_N0
cycloneive_ram_block ram_block3a23(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a23_PORTADATAOUT_bus),
	.portbdataout(ram_block3a23_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a23.clk0_core_clock_enable = "ena0";
defparam ram_block3a23.clk1_core_clock_enable = "ena1";
defparam ram_block3a23.data_interleave_offset_in_bits = 1;
defparam ram_block3a23.data_interleave_width_in_bits = 1;
defparam ram_block3a23.init_file = "meminit.hex";
defparam ram_block3a23.init_file_layout = "port_a";
defparam ram_block3a23.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a23.operation_mode = "bidir_dual_port";
defparam ram_block3a23.port_a_address_clear = "none";
defparam ram_block3a23.port_a_address_width = 13;
defparam ram_block3a23.port_a_byte_enable_clock = "none";
defparam ram_block3a23.port_a_data_out_clear = "none";
defparam ram_block3a23.port_a_data_out_clock = "none";
defparam ram_block3a23.port_a_data_width = 1;
defparam ram_block3a23.port_a_first_address = 0;
defparam ram_block3a23.port_a_first_bit_number = 23;
defparam ram_block3a23.port_a_last_address = 8191;
defparam ram_block3a23.port_a_logical_ram_depth = 16384;
defparam ram_block3a23.port_a_logical_ram_width = 32;
defparam ram_block3a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_address_clear = "none";
defparam ram_block3a23.port_b_address_clock = "clock1";
defparam ram_block3a23.port_b_address_width = 13;
defparam ram_block3a23.port_b_data_in_clock = "clock1";
defparam ram_block3a23.port_b_data_out_clear = "none";
defparam ram_block3a23.port_b_data_out_clock = "none";
defparam ram_block3a23.port_b_data_width = 1;
defparam ram_block3a23.port_b_first_address = 0;
defparam ram_block3a23.port_b_first_bit_number = 23;
defparam ram_block3a23.port_b_last_address = 8191;
defparam ram_block3a23.port_b_logical_ram_depth = 16384;
defparam ram_block3a23.port_b_logical_ram_width = 32;
defparam ram_block3a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_read_enable_clock = "clock1";
defparam ram_block3a23.port_b_write_enable_clock = "clock1";
defparam ram_block3a23.ram_block_type = "M9K";
defparam ram_block3a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E5CB187BC004B601000;
// synopsys translate_on

// Location: M9K_X64_Y36_N0
cycloneive_ram_block ram_block3a56(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a56_PORTADATAOUT_bus),
	.portbdataout(ram_block3a56_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a56.clk0_core_clock_enable = "ena0";
defparam ram_block3a56.clk1_core_clock_enable = "ena1";
defparam ram_block3a56.data_interleave_offset_in_bits = 1;
defparam ram_block3a56.data_interleave_width_in_bits = 1;
defparam ram_block3a56.init_file = "meminit.hex";
defparam ram_block3a56.init_file_layout = "port_a";
defparam ram_block3a56.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a56.operation_mode = "bidir_dual_port";
defparam ram_block3a56.port_a_address_clear = "none";
defparam ram_block3a56.port_a_address_width = 13;
defparam ram_block3a56.port_a_byte_enable_clock = "none";
defparam ram_block3a56.port_a_data_out_clear = "none";
defparam ram_block3a56.port_a_data_out_clock = "none";
defparam ram_block3a56.port_a_data_width = 1;
defparam ram_block3a56.port_a_first_address = 0;
defparam ram_block3a56.port_a_first_bit_number = 24;
defparam ram_block3a56.port_a_last_address = 8191;
defparam ram_block3a56.port_a_logical_ram_depth = 16384;
defparam ram_block3a56.port_a_logical_ram_width = 32;
defparam ram_block3a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_address_clear = "none";
defparam ram_block3a56.port_b_address_clock = "clock1";
defparam ram_block3a56.port_b_address_width = 13;
defparam ram_block3a56.port_b_data_in_clock = "clock1";
defparam ram_block3a56.port_b_data_out_clear = "none";
defparam ram_block3a56.port_b_data_out_clock = "none";
defparam ram_block3a56.port_b_data_width = 1;
defparam ram_block3a56.port_b_first_address = 0;
defparam ram_block3a56.port_b_first_bit_number = 24;
defparam ram_block3a56.port_b_last_address = 8191;
defparam ram_block3a56.port_b_logical_ram_depth = 16384;
defparam ram_block3a56.port_b_logical_ram_width = 32;
defparam ram_block3a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_read_enable_clock = "clock1";
defparam ram_block3a56.port_b_write_enable_clock = "clock1";
defparam ram_block3a56.ram_block_type = "M9K";
defparam ram_block3a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y41_N0
cycloneive_ram_block ram_block3a24(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a24_PORTADATAOUT_bus),
	.portbdataout(ram_block3a24_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a24.clk0_core_clock_enable = "ena0";
defparam ram_block3a24.clk1_core_clock_enable = "ena1";
defparam ram_block3a24.data_interleave_offset_in_bits = 1;
defparam ram_block3a24.data_interleave_width_in_bits = 1;
defparam ram_block3a24.init_file = "meminit.hex";
defparam ram_block3a24.init_file_layout = "port_a";
defparam ram_block3a24.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a24.operation_mode = "bidir_dual_port";
defparam ram_block3a24.port_a_address_clear = "none";
defparam ram_block3a24.port_a_address_width = 13;
defparam ram_block3a24.port_a_byte_enable_clock = "none";
defparam ram_block3a24.port_a_data_out_clear = "none";
defparam ram_block3a24.port_a_data_out_clock = "none";
defparam ram_block3a24.port_a_data_width = 1;
defparam ram_block3a24.port_a_first_address = 0;
defparam ram_block3a24.port_a_first_bit_number = 24;
defparam ram_block3a24.port_a_last_address = 8191;
defparam ram_block3a24.port_a_logical_ram_depth = 16384;
defparam ram_block3a24.port_a_logical_ram_width = 32;
defparam ram_block3a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_address_clear = "none";
defparam ram_block3a24.port_b_address_clock = "clock1";
defparam ram_block3a24.port_b_address_width = 13;
defparam ram_block3a24.port_b_data_in_clock = "clock1";
defparam ram_block3a24.port_b_data_out_clear = "none";
defparam ram_block3a24.port_b_data_out_clock = "none";
defparam ram_block3a24.port_b_data_width = 1;
defparam ram_block3a24.port_b_first_address = 0;
defparam ram_block3a24.port_b_first_bit_number = 24;
defparam ram_block3a24.port_b_last_address = 8191;
defparam ram_block3a24.port_b_logical_ram_depth = 16384;
defparam ram_block3a24.port_b_logical_ram_width = 32;
defparam ram_block3a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_read_enable_clock = "clock1";
defparam ram_block3a24.port_b_write_enable_clock = "clock1";
defparam ram_block3a24.ram_block_type = "M9K";
defparam ram_block3a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021830C680DB793600400;
// synopsys translate_on

// Location: M9K_X37_Y32_N0
cycloneive_ram_block ram_block3a57(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a57_PORTADATAOUT_bus),
	.portbdataout(ram_block3a57_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a57.clk0_core_clock_enable = "ena0";
defparam ram_block3a57.clk1_core_clock_enable = "ena1";
defparam ram_block3a57.data_interleave_offset_in_bits = 1;
defparam ram_block3a57.data_interleave_width_in_bits = 1;
defparam ram_block3a57.init_file = "meminit.hex";
defparam ram_block3a57.init_file_layout = "port_a";
defparam ram_block3a57.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a57.operation_mode = "bidir_dual_port";
defparam ram_block3a57.port_a_address_clear = "none";
defparam ram_block3a57.port_a_address_width = 13;
defparam ram_block3a57.port_a_byte_enable_clock = "none";
defparam ram_block3a57.port_a_data_out_clear = "none";
defparam ram_block3a57.port_a_data_out_clock = "none";
defparam ram_block3a57.port_a_data_width = 1;
defparam ram_block3a57.port_a_first_address = 0;
defparam ram_block3a57.port_a_first_bit_number = 25;
defparam ram_block3a57.port_a_last_address = 8191;
defparam ram_block3a57.port_a_logical_ram_depth = 16384;
defparam ram_block3a57.port_a_logical_ram_width = 32;
defparam ram_block3a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_address_clear = "none";
defparam ram_block3a57.port_b_address_clock = "clock1";
defparam ram_block3a57.port_b_address_width = 13;
defparam ram_block3a57.port_b_data_in_clock = "clock1";
defparam ram_block3a57.port_b_data_out_clear = "none";
defparam ram_block3a57.port_b_data_out_clock = "none";
defparam ram_block3a57.port_b_data_width = 1;
defparam ram_block3a57.port_b_first_address = 0;
defparam ram_block3a57.port_b_first_bit_number = 25;
defparam ram_block3a57.port_b_last_address = 8191;
defparam ram_block3a57.port_b_logical_ram_depth = 16384;
defparam ram_block3a57.port_b_logical_ram_width = 32;
defparam ram_block3a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_read_enable_clock = "clock1";
defparam ram_block3a57.port_b_write_enable_clock = "clock1";
defparam ram_block3a57.ram_block_type = "M9K";
defparam ram_block3a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y48_N0
cycloneive_ram_block ram_block3a25(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a25_PORTADATAOUT_bus),
	.portbdataout(ram_block3a25_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a25.clk0_core_clock_enable = "ena0";
defparam ram_block3a25.clk1_core_clock_enable = "ena1";
defparam ram_block3a25.data_interleave_offset_in_bits = 1;
defparam ram_block3a25.data_interleave_width_in_bits = 1;
defparam ram_block3a25.init_file = "meminit.hex";
defparam ram_block3a25.init_file_layout = "port_a";
defparam ram_block3a25.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a25.operation_mode = "bidir_dual_port";
defparam ram_block3a25.port_a_address_clear = "none";
defparam ram_block3a25.port_a_address_width = 13;
defparam ram_block3a25.port_a_byte_enable_clock = "none";
defparam ram_block3a25.port_a_data_out_clear = "none";
defparam ram_block3a25.port_a_data_out_clock = "none";
defparam ram_block3a25.port_a_data_width = 1;
defparam ram_block3a25.port_a_first_address = 0;
defparam ram_block3a25.port_a_first_bit_number = 25;
defparam ram_block3a25.port_a_last_address = 8191;
defparam ram_block3a25.port_a_logical_ram_depth = 16384;
defparam ram_block3a25.port_a_logical_ram_width = 32;
defparam ram_block3a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_address_clear = "none";
defparam ram_block3a25.port_b_address_clock = "clock1";
defparam ram_block3a25.port_b_address_width = 13;
defparam ram_block3a25.port_b_data_in_clock = "clock1";
defparam ram_block3a25.port_b_data_out_clear = "none";
defparam ram_block3a25.port_b_data_out_clock = "none";
defparam ram_block3a25.port_b_data_width = 1;
defparam ram_block3a25.port_b_first_address = 0;
defparam ram_block3a25.port_b_first_bit_number = 25;
defparam ram_block3a25.port_b_last_address = 8191;
defparam ram_block3a25.port_b_logical_ram_depth = 16384;
defparam ram_block3a25.port_b_logical_ram_width = 32;
defparam ram_block3a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_read_enable_clock = "clock1";
defparam ram_block3a25.port_b_write_enable_clock = "clock1";
defparam ram_block3a25.ram_block_type = "M9K";
defparam ram_block3a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000CB783600310;
// synopsys translate_on

// Location: M9K_X78_Y38_N0
cycloneive_ram_block ram_block3a58(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a58_PORTADATAOUT_bus),
	.portbdataout(ram_block3a58_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a58.clk0_core_clock_enable = "ena0";
defparam ram_block3a58.clk1_core_clock_enable = "ena1";
defparam ram_block3a58.data_interleave_offset_in_bits = 1;
defparam ram_block3a58.data_interleave_width_in_bits = 1;
defparam ram_block3a58.init_file = "meminit.hex";
defparam ram_block3a58.init_file_layout = "port_a";
defparam ram_block3a58.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a58.operation_mode = "bidir_dual_port";
defparam ram_block3a58.port_a_address_clear = "none";
defparam ram_block3a58.port_a_address_width = 13;
defparam ram_block3a58.port_a_byte_enable_clock = "none";
defparam ram_block3a58.port_a_data_out_clear = "none";
defparam ram_block3a58.port_a_data_out_clock = "none";
defparam ram_block3a58.port_a_data_width = 1;
defparam ram_block3a58.port_a_first_address = 0;
defparam ram_block3a58.port_a_first_bit_number = 26;
defparam ram_block3a58.port_a_last_address = 8191;
defparam ram_block3a58.port_a_logical_ram_depth = 16384;
defparam ram_block3a58.port_a_logical_ram_width = 32;
defparam ram_block3a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_address_clear = "none";
defparam ram_block3a58.port_b_address_clock = "clock1";
defparam ram_block3a58.port_b_address_width = 13;
defparam ram_block3a58.port_b_data_in_clock = "clock1";
defparam ram_block3a58.port_b_data_out_clear = "none";
defparam ram_block3a58.port_b_data_out_clock = "none";
defparam ram_block3a58.port_b_data_width = 1;
defparam ram_block3a58.port_b_first_address = 0;
defparam ram_block3a58.port_b_first_bit_number = 26;
defparam ram_block3a58.port_b_last_address = 8191;
defparam ram_block3a58.port_b_logical_ram_depth = 16384;
defparam ram_block3a58.port_b_logical_ram_width = 32;
defparam ram_block3a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_read_enable_clock = "clock1";
defparam ram_block3a58.port_b_write_enable_clock = "clock1";
defparam ram_block3a58.ram_block_type = "M9K";
defparam ram_block3a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y39_N0
cycloneive_ram_block ram_block3a26(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a26_PORTADATAOUT_bus),
	.portbdataout(ram_block3a26_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a26.clk0_core_clock_enable = "ena0";
defparam ram_block3a26.clk1_core_clock_enable = "ena1";
defparam ram_block3a26.data_interleave_offset_in_bits = 1;
defparam ram_block3a26.data_interleave_width_in_bits = 1;
defparam ram_block3a26.init_file = "meminit.hex";
defparam ram_block3a26.init_file_layout = "port_a";
defparam ram_block3a26.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a26.operation_mode = "bidir_dual_port";
defparam ram_block3a26.port_a_address_clear = "none";
defparam ram_block3a26.port_a_address_width = 13;
defparam ram_block3a26.port_a_byte_enable_clock = "none";
defparam ram_block3a26.port_a_data_out_clear = "none";
defparam ram_block3a26.port_a_data_out_clock = "none";
defparam ram_block3a26.port_a_data_width = 1;
defparam ram_block3a26.port_a_first_address = 0;
defparam ram_block3a26.port_a_first_bit_number = 26;
defparam ram_block3a26.port_a_last_address = 8191;
defparam ram_block3a26.port_a_logical_ram_depth = 16384;
defparam ram_block3a26.port_a_logical_ram_width = 32;
defparam ram_block3a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_address_clear = "none";
defparam ram_block3a26.port_b_address_clock = "clock1";
defparam ram_block3a26.port_b_address_width = 13;
defparam ram_block3a26.port_b_data_in_clock = "clock1";
defparam ram_block3a26.port_b_data_out_clear = "none";
defparam ram_block3a26.port_b_data_out_clock = "none";
defparam ram_block3a26.port_b_data_width = 1;
defparam ram_block3a26.port_b_first_address = 0;
defparam ram_block3a26.port_b_first_bit_number = 26;
defparam ram_block3a26.port_b_last_address = 8191;
defparam ram_block3a26.port_b_logical_ram_depth = 16384;
defparam ram_block3a26.port_b_logical_ram_width = 32;
defparam ram_block3a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_read_enable_clock = "clock1";
defparam ram_block3a26.port_b_write_enable_clock = "clock1";
defparam ram_block3a26.ram_block_type = "M9K";
defparam ram_block3a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007CFBDE639B287F0888F;
// synopsys translate_on

// Location: M9K_X51_Y46_N0
cycloneive_ram_block ram_block3a59(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a59_PORTADATAOUT_bus),
	.portbdataout(ram_block3a59_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a59.clk0_core_clock_enable = "ena0";
defparam ram_block3a59.clk1_core_clock_enable = "ena1";
defparam ram_block3a59.data_interleave_offset_in_bits = 1;
defparam ram_block3a59.data_interleave_width_in_bits = 1;
defparam ram_block3a59.init_file = "meminit.hex";
defparam ram_block3a59.init_file_layout = "port_a";
defparam ram_block3a59.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a59.operation_mode = "bidir_dual_port";
defparam ram_block3a59.port_a_address_clear = "none";
defparam ram_block3a59.port_a_address_width = 13;
defparam ram_block3a59.port_a_byte_enable_clock = "none";
defparam ram_block3a59.port_a_data_out_clear = "none";
defparam ram_block3a59.port_a_data_out_clock = "none";
defparam ram_block3a59.port_a_data_width = 1;
defparam ram_block3a59.port_a_first_address = 0;
defparam ram_block3a59.port_a_first_bit_number = 27;
defparam ram_block3a59.port_a_last_address = 8191;
defparam ram_block3a59.port_a_logical_ram_depth = 16384;
defparam ram_block3a59.port_a_logical_ram_width = 32;
defparam ram_block3a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_address_clear = "none";
defparam ram_block3a59.port_b_address_clock = "clock1";
defparam ram_block3a59.port_b_address_width = 13;
defparam ram_block3a59.port_b_data_in_clock = "clock1";
defparam ram_block3a59.port_b_data_out_clear = "none";
defparam ram_block3a59.port_b_data_out_clock = "none";
defparam ram_block3a59.port_b_data_width = 1;
defparam ram_block3a59.port_b_first_address = 0;
defparam ram_block3a59.port_b_first_bit_number = 27;
defparam ram_block3a59.port_b_last_address = 8191;
defparam ram_block3a59.port_b_logical_ram_depth = 16384;
defparam ram_block3a59.port_b_logical_ram_width = 32;
defparam ram_block3a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_read_enable_clock = "clock1";
defparam ram_block3a59.port_b_write_enable_clock = "clock1";
defparam ram_block3a59.ram_block_type = "M9K";
defparam ram_block3a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y32_N0
cycloneive_ram_block ram_block3a27(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a27_PORTADATAOUT_bus),
	.portbdataout(ram_block3a27_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a27.clk0_core_clock_enable = "ena0";
defparam ram_block3a27.clk1_core_clock_enable = "ena1";
defparam ram_block3a27.data_interleave_offset_in_bits = 1;
defparam ram_block3a27.data_interleave_width_in_bits = 1;
defparam ram_block3a27.init_file = "meminit.hex";
defparam ram_block3a27.init_file_layout = "port_a";
defparam ram_block3a27.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a27.operation_mode = "bidir_dual_port";
defparam ram_block3a27.port_a_address_clear = "none";
defparam ram_block3a27.port_a_address_width = 13;
defparam ram_block3a27.port_a_byte_enable_clock = "none";
defparam ram_block3a27.port_a_data_out_clear = "none";
defparam ram_block3a27.port_a_data_out_clock = "none";
defparam ram_block3a27.port_a_data_width = 1;
defparam ram_block3a27.port_a_first_address = 0;
defparam ram_block3a27.port_a_first_bit_number = 27;
defparam ram_block3a27.port_a_last_address = 8191;
defparam ram_block3a27.port_a_logical_ram_depth = 16384;
defparam ram_block3a27.port_a_logical_ram_width = 32;
defparam ram_block3a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_address_clear = "none";
defparam ram_block3a27.port_b_address_clock = "clock1";
defparam ram_block3a27.port_b_address_width = 13;
defparam ram_block3a27.port_b_data_in_clock = "clock1";
defparam ram_block3a27.port_b_data_out_clear = "none";
defparam ram_block3a27.port_b_data_out_clock = "none";
defparam ram_block3a27.port_b_data_width = 1;
defparam ram_block3a27.port_b_first_address = 0;
defparam ram_block3a27.port_b_first_bit_number = 27;
defparam ram_block3a27.port_b_last_address = 8191;
defparam ram_block3a27.port_b_logical_ram_depth = 16384;
defparam ram_block3a27.port_b_logical_ram_width = 32;
defparam ram_block3a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_read_enable_clock = "clock1";
defparam ram_block3a27.port_b_write_enable_clock = "clock1";
defparam ram_block3a27.ram_block_type = "M9K";
defparam ram_block3a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010E1C6264AD282C08088;
// synopsys translate_on

// Location: M9K_X51_Y38_N0
cycloneive_ram_block ram_block3a60(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a60_PORTADATAOUT_bus),
	.portbdataout(ram_block3a60_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a60.clk0_core_clock_enable = "ena0";
defparam ram_block3a60.clk1_core_clock_enable = "ena1";
defparam ram_block3a60.data_interleave_offset_in_bits = 1;
defparam ram_block3a60.data_interleave_width_in_bits = 1;
defparam ram_block3a60.init_file = "meminit.hex";
defparam ram_block3a60.init_file_layout = "port_a";
defparam ram_block3a60.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a60.operation_mode = "bidir_dual_port";
defparam ram_block3a60.port_a_address_clear = "none";
defparam ram_block3a60.port_a_address_width = 13;
defparam ram_block3a60.port_a_byte_enable_clock = "none";
defparam ram_block3a60.port_a_data_out_clear = "none";
defparam ram_block3a60.port_a_data_out_clock = "none";
defparam ram_block3a60.port_a_data_width = 1;
defparam ram_block3a60.port_a_first_address = 0;
defparam ram_block3a60.port_a_first_bit_number = 28;
defparam ram_block3a60.port_a_last_address = 8191;
defparam ram_block3a60.port_a_logical_ram_depth = 16384;
defparam ram_block3a60.port_a_logical_ram_width = 32;
defparam ram_block3a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_address_clear = "none";
defparam ram_block3a60.port_b_address_clock = "clock1";
defparam ram_block3a60.port_b_address_width = 13;
defparam ram_block3a60.port_b_data_in_clock = "clock1";
defparam ram_block3a60.port_b_data_out_clear = "none";
defparam ram_block3a60.port_b_data_out_clock = "none";
defparam ram_block3a60.port_b_data_width = 1;
defparam ram_block3a60.port_b_first_address = 0;
defparam ram_block3a60.port_b_first_bit_number = 28;
defparam ram_block3a60.port_b_last_address = 8191;
defparam ram_block3a60.port_b_logical_ram_depth = 16384;
defparam ram_block3a60.port_b_logical_ram_width = 32;
defparam ram_block3a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_read_enable_clock = "clock1";
defparam ram_block3a60.port_b_write_enable_clock = "clock1";
defparam ram_block3a60.ram_block_type = "M9K";
defparam ram_block3a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y40_N0
cycloneive_ram_block ram_block3a28(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a28_PORTADATAOUT_bus),
	.portbdataout(ram_block3a28_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a28.clk0_core_clock_enable = "ena0";
defparam ram_block3a28.clk1_core_clock_enable = "ena1";
defparam ram_block3a28.data_interleave_offset_in_bits = 1;
defparam ram_block3a28.data_interleave_width_in_bits = 1;
defparam ram_block3a28.init_file = "meminit.hex";
defparam ram_block3a28.init_file_layout = "port_a";
defparam ram_block3a28.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a28.operation_mode = "bidir_dual_port";
defparam ram_block3a28.port_a_address_clear = "none";
defparam ram_block3a28.port_a_address_width = 13;
defparam ram_block3a28.port_a_byte_enable_clock = "none";
defparam ram_block3a28.port_a_data_out_clear = "none";
defparam ram_block3a28.port_a_data_out_clock = "none";
defparam ram_block3a28.port_a_data_width = 1;
defparam ram_block3a28.port_a_first_address = 0;
defparam ram_block3a28.port_a_first_bit_number = 28;
defparam ram_block3a28.port_a_last_address = 8191;
defparam ram_block3a28.port_a_logical_ram_depth = 16384;
defparam ram_block3a28.port_a_logical_ram_width = 32;
defparam ram_block3a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_address_clear = "none";
defparam ram_block3a28.port_b_address_clock = "clock1";
defparam ram_block3a28.port_b_address_width = 13;
defparam ram_block3a28.port_b_data_in_clock = "clock1";
defparam ram_block3a28.port_b_data_out_clear = "none";
defparam ram_block3a28.port_b_data_out_clock = "none";
defparam ram_block3a28.port_b_data_width = 1;
defparam ram_block3a28.port_b_first_address = 0;
defparam ram_block3a28.port_b_first_bit_number = 28;
defparam ram_block3a28.port_b_last_address = 8191;
defparam ram_block3a28.port_b_logical_ram_depth = 16384;
defparam ram_block3a28.port_b_logical_ram_width = 32;
defparam ram_block3a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_read_enable_clock = "clock1";
defparam ram_block3a28.port_b_write_enable_clock = "clock1";
defparam ram_block3a28.ram_block_type = "M9K";
defparam ram_block3a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008100011B00926100807;
// synopsys translate_on

// Location: M9K_X64_Y39_N0
cycloneive_ram_block ram_block3a61(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a61_PORTADATAOUT_bus),
	.portbdataout(ram_block3a61_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a61.clk0_core_clock_enable = "ena0";
defparam ram_block3a61.clk1_core_clock_enable = "ena1";
defparam ram_block3a61.data_interleave_offset_in_bits = 1;
defparam ram_block3a61.data_interleave_width_in_bits = 1;
defparam ram_block3a61.init_file = "meminit.hex";
defparam ram_block3a61.init_file_layout = "port_a";
defparam ram_block3a61.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a61.operation_mode = "bidir_dual_port";
defparam ram_block3a61.port_a_address_clear = "none";
defparam ram_block3a61.port_a_address_width = 13;
defparam ram_block3a61.port_a_byte_enable_clock = "none";
defparam ram_block3a61.port_a_data_out_clear = "none";
defparam ram_block3a61.port_a_data_out_clock = "none";
defparam ram_block3a61.port_a_data_width = 1;
defparam ram_block3a61.port_a_first_address = 0;
defparam ram_block3a61.port_a_first_bit_number = 29;
defparam ram_block3a61.port_a_last_address = 8191;
defparam ram_block3a61.port_a_logical_ram_depth = 16384;
defparam ram_block3a61.port_a_logical_ram_width = 32;
defparam ram_block3a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_address_clear = "none";
defparam ram_block3a61.port_b_address_clock = "clock1";
defparam ram_block3a61.port_b_address_width = 13;
defparam ram_block3a61.port_b_data_in_clock = "clock1";
defparam ram_block3a61.port_b_data_out_clear = "none";
defparam ram_block3a61.port_b_data_out_clock = "none";
defparam ram_block3a61.port_b_data_width = 1;
defparam ram_block3a61.port_b_first_address = 0;
defparam ram_block3a61.port_b_first_bit_number = 29;
defparam ram_block3a61.port_b_last_address = 8191;
defparam ram_block3a61.port_b_logical_ram_depth = 16384;
defparam ram_block3a61.port_b_logical_ram_width = 32;
defparam ram_block3a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_read_enable_clock = "clock1";
defparam ram_block3a61.port_b_write_enable_clock = "clock1";
defparam ram_block3a61.ram_block_type = "M9K";
defparam ram_block3a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y39_N0
cycloneive_ram_block ram_block3a29(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a29_PORTADATAOUT_bus),
	.portbdataout(ram_block3a29_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a29.clk0_core_clock_enable = "ena0";
defparam ram_block3a29.clk1_core_clock_enable = "ena1";
defparam ram_block3a29.data_interleave_offset_in_bits = 1;
defparam ram_block3a29.data_interleave_width_in_bits = 1;
defparam ram_block3a29.init_file = "meminit.hex";
defparam ram_block3a29.init_file_layout = "port_a";
defparam ram_block3a29.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a29.operation_mode = "bidir_dual_port";
defparam ram_block3a29.port_a_address_clear = "none";
defparam ram_block3a29.port_a_address_width = 13;
defparam ram_block3a29.port_a_byte_enable_clock = "none";
defparam ram_block3a29.port_a_data_out_clear = "none";
defparam ram_block3a29.port_a_data_out_clock = "none";
defparam ram_block3a29.port_a_data_width = 1;
defparam ram_block3a29.port_a_first_address = 0;
defparam ram_block3a29.port_a_first_bit_number = 29;
defparam ram_block3a29.port_a_last_address = 8191;
defparam ram_block3a29.port_a_logical_ram_depth = 16384;
defparam ram_block3a29.port_a_logical_ram_width = 32;
defparam ram_block3a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_address_clear = "none";
defparam ram_block3a29.port_b_address_clock = "clock1";
defparam ram_block3a29.port_b_address_width = 13;
defparam ram_block3a29.port_b_data_in_clock = "clock1";
defparam ram_block3a29.port_b_data_out_clear = "none";
defparam ram_block3a29.port_b_data_out_clock = "none";
defparam ram_block3a29.port_b_data_width = 1;
defparam ram_block3a29.port_b_first_address = 0;
defparam ram_block3a29.port_b_first_bit_number = 29;
defparam ram_block3a29.port_b_last_address = 8191;
defparam ram_block3a29.port_b_logical_ram_depth = 16384;
defparam ram_block3a29.port_b_logical_ram_width = 32;
defparam ram_block3a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_read_enable_clock = "clock1";
defparam ram_block3a29.port_b_write_enable_clock = "clock1";
defparam ram_block3a29.ram_block_type = "M9K";
defparam ram_block3a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000078F3DE001B007700807;
// synopsys translate_on

// Location: M9K_X78_Y42_N0
cycloneive_ram_block ram_block3a62(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a62_PORTADATAOUT_bus),
	.portbdataout(ram_block3a62_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a62.clk0_core_clock_enable = "ena0";
defparam ram_block3a62.clk1_core_clock_enable = "ena1";
defparam ram_block3a62.data_interleave_offset_in_bits = 1;
defparam ram_block3a62.data_interleave_width_in_bits = 1;
defparam ram_block3a62.init_file = "meminit.hex";
defparam ram_block3a62.init_file_layout = "port_a";
defparam ram_block3a62.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a62.operation_mode = "bidir_dual_port";
defparam ram_block3a62.port_a_address_clear = "none";
defparam ram_block3a62.port_a_address_width = 13;
defparam ram_block3a62.port_a_byte_enable_clock = "none";
defparam ram_block3a62.port_a_data_out_clear = "none";
defparam ram_block3a62.port_a_data_out_clock = "none";
defparam ram_block3a62.port_a_data_width = 1;
defparam ram_block3a62.port_a_first_address = 0;
defparam ram_block3a62.port_a_first_bit_number = 30;
defparam ram_block3a62.port_a_last_address = 8191;
defparam ram_block3a62.port_a_logical_ram_depth = 16384;
defparam ram_block3a62.port_a_logical_ram_width = 32;
defparam ram_block3a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_address_clear = "none";
defparam ram_block3a62.port_b_address_clock = "clock1";
defparam ram_block3a62.port_b_address_width = 13;
defparam ram_block3a62.port_b_data_in_clock = "clock1";
defparam ram_block3a62.port_b_data_out_clear = "none";
defparam ram_block3a62.port_b_data_out_clock = "none";
defparam ram_block3a62.port_b_data_width = 1;
defparam ram_block3a62.port_b_first_address = 0;
defparam ram_block3a62.port_b_first_bit_number = 30;
defparam ram_block3a62.port_b_last_address = 8191;
defparam ram_block3a62.port_b_logical_ram_depth = 16384;
defparam ram_block3a62.port_b_logical_ram_width = 32;
defparam ram_block3a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_read_enable_clock = "clock1";
defparam ram_block3a62.port_b_write_enable_clock = "clock1";
defparam ram_block3a62.ram_block_type = "M9K";
defparam ram_block3a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y42_N0
cycloneive_ram_block ram_block3a30(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a30_PORTADATAOUT_bus),
	.portbdataout(ram_block3a30_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a30.clk0_core_clock_enable = "ena0";
defparam ram_block3a30.clk1_core_clock_enable = "ena1";
defparam ram_block3a30.data_interleave_offset_in_bits = 1;
defparam ram_block3a30.data_interleave_width_in_bits = 1;
defparam ram_block3a30.init_file = "meminit.hex";
defparam ram_block3a30.init_file_layout = "port_a";
defparam ram_block3a30.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a30.operation_mode = "bidir_dual_port";
defparam ram_block3a30.port_a_address_clear = "none";
defparam ram_block3a30.port_a_address_width = 13;
defparam ram_block3a30.port_a_byte_enable_clock = "none";
defparam ram_block3a30.port_a_data_out_clear = "none";
defparam ram_block3a30.port_a_data_out_clock = "none";
defparam ram_block3a30.port_a_data_width = 1;
defparam ram_block3a30.port_a_first_address = 0;
defparam ram_block3a30.port_a_first_bit_number = 30;
defparam ram_block3a30.port_a_last_address = 8191;
defparam ram_block3a30.port_a_logical_ram_depth = 16384;
defparam ram_block3a30.port_a_logical_ram_width = 32;
defparam ram_block3a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_address_clear = "none";
defparam ram_block3a30.port_b_address_clock = "clock1";
defparam ram_block3a30.port_b_address_width = 13;
defparam ram_block3a30.port_b_data_in_clock = "clock1";
defparam ram_block3a30.port_b_data_out_clear = "none";
defparam ram_block3a30.port_b_data_out_clock = "none";
defparam ram_block3a30.port_b_data_width = 1;
defparam ram_block3a30.port_b_first_address = 0;
defparam ram_block3a30.port_b_first_bit_number = 30;
defparam ram_block3a30.port_b_last_address = 8191;
defparam ram_block3a30.port_b_logical_ram_depth = 16384;
defparam ram_block3a30.port_b_logical_ram_width = 32;
defparam ram_block3a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_read_enable_clock = "clock1";
defparam ram_block3a30.port_b_write_enable_clock = "clock1";
defparam ram_block3a30.ram_block_type = "M9K";
defparam ram_block3a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000;
// synopsys translate_on

// Location: M9K_X37_Y40_N0
cycloneive_ram_block ram_block3a63(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a63_PORTADATAOUT_bus),
	.portbdataout(ram_block3a63_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a63.clk0_core_clock_enable = "ena0";
defparam ram_block3a63.clk1_core_clock_enable = "ena1";
defparam ram_block3a63.data_interleave_offset_in_bits = 1;
defparam ram_block3a63.data_interleave_width_in_bits = 1;
defparam ram_block3a63.init_file = "meminit.hex";
defparam ram_block3a63.init_file_layout = "port_a";
defparam ram_block3a63.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a63.operation_mode = "bidir_dual_port";
defparam ram_block3a63.port_a_address_clear = "none";
defparam ram_block3a63.port_a_address_width = 13;
defparam ram_block3a63.port_a_byte_enable_clock = "none";
defparam ram_block3a63.port_a_data_out_clear = "none";
defparam ram_block3a63.port_a_data_out_clock = "none";
defparam ram_block3a63.port_a_data_width = 1;
defparam ram_block3a63.port_a_first_address = 0;
defparam ram_block3a63.port_a_first_bit_number = 31;
defparam ram_block3a63.port_a_last_address = 8191;
defparam ram_block3a63.port_a_logical_ram_depth = 16384;
defparam ram_block3a63.port_a_logical_ram_width = 32;
defparam ram_block3a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_address_clear = "none";
defparam ram_block3a63.port_b_address_clock = "clock1";
defparam ram_block3a63.port_b_address_width = 13;
defparam ram_block3a63.port_b_data_in_clock = "clock1";
defparam ram_block3a63.port_b_data_out_clear = "none";
defparam ram_block3a63.port_b_data_out_clock = "none";
defparam ram_block3a63.port_b_data_width = 1;
defparam ram_block3a63.port_b_first_address = 0;
defparam ram_block3a63.port_b_first_bit_number = 31;
defparam ram_block3a63.port_b_last_address = 8191;
defparam ram_block3a63.port_b_logical_ram_depth = 16384;
defparam ram_block3a63.port_b_logical_ram_width = 32;
defparam ram_block3a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_read_enable_clock = "clock1";
defparam ram_block3a63.port_b_write_enable_clock = "clock1";
defparam ram_block3a63.ram_block_type = "M9K";
defparam ram_block3a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y40_N0
cycloneive_ram_block ram_block3a31(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a31_PORTADATAOUT_bus),
	.portbdataout(ram_block3a31_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a31.clk0_core_clock_enable = "ena0";
defparam ram_block3a31.clk1_core_clock_enable = "ena1";
defparam ram_block3a31.data_interleave_offset_in_bits = 1;
defparam ram_block3a31.data_interleave_width_in_bits = 1;
defparam ram_block3a31.init_file = "meminit.hex";
defparam ram_block3a31.init_file_layout = "port_a";
defparam ram_block3a31.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a31.operation_mode = "bidir_dual_port";
defparam ram_block3a31.port_a_address_clear = "none";
defparam ram_block3a31.port_a_address_width = 13;
defparam ram_block3a31.port_a_byte_enable_clock = "none";
defparam ram_block3a31.port_a_data_out_clear = "none";
defparam ram_block3a31.port_a_data_out_clock = "none";
defparam ram_block3a31.port_a_data_width = 1;
defparam ram_block3a31.port_a_first_address = 0;
defparam ram_block3a31.port_a_first_bit_number = 31;
defparam ram_block3a31.port_a_last_address = 8191;
defparam ram_block3a31.port_a_logical_ram_depth = 16384;
defparam ram_block3a31.port_a_logical_ram_width = 32;
defparam ram_block3a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_address_clear = "none";
defparam ram_block3a31.port_b_address_clock = "clock1";
defparam ram_block3a31.port_b_address_width = 13;
defparam ram_block3a31.port_b_data_in_clock = "clock1";
defparam ram_block3a31.port_b_data_out_clear = "none";
defparam ram_block3a31.port_b_data_out_clock = "none";
defparam ram_block3a31.port_b_data_width = 1;
defparam ram_block3a31.port_b_first_address = 0;
defparam ram_block3a31.port_b_first_bit_number = 31;
defparam ram_block3a31.port_b_last_address = 8191;
defparam ram_block3a31.port_b_logical_ram_depth = 16384;
defparam ram_block3a31.port_b_logical_ram_width = 32;
defparam ram_block3a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_read_enable_clock = "clock1";
defparam ram_block3a31.port_b_write_enable_clock = "clock1";
defparam ram_block3a31.ram_block_type = "M9K";
defparam ram_block3a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000C18426089282400008;
// synopsys translate_on

// Location: FF_X55_Y37_N29
dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_a_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N31
dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(\address_reg_b[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_b_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N30
cycloneive_lcell_comb \address_reg_b[0]~feeder (
// Equation(s):
// \address_reg_b[0]~feeder_combout  = ram_rom_addr_reg_13

	.dataa(gnd),
	.datab(gnd),
	.datac(ram_rom_addr_reg_13),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg_b[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_b[0]~feeder .lut_mask = 16'hF0F0;
defparam \address_reg_b[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa (
	ramaddr,
	ramWEN,
	always1,
	eq_node_1,
	eq_node_0,
	devpor,
	devclrn,
	devoe);
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	eq_node_1;
output 	eq_node_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X59_Y34_N28
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (!\ramWEN~0_combout  & (!\ramaddr~29_combout  & always1))

	.dataa(ramWEN),
	.datab(gnd),
	.datac(ramaddr),
	.datad(always1),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h0500;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N2
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (!\ramWEN~0_combout  & (always1 & \ramaddr~29_combout ))

	.dataa(ramWEN),
	.datab(always1),
	.datac(gnd),
	.datad(ramaddr),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h4400;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa_1 (
	ram_rom_addr_reg_13,
	sdr,
	eq_node_1,
	eq_node_0,
	irf_reg_2_1,
	state_5,
	devpor,
	devclrn,
	devoe);
input 	ram_rom_addr_reg_13;
input 	sdr;
output 	eq_node_1;
output 	eq_node_0;
input 	irf_reg_2_1;
input 	state_5;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X48_Y37_N24
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (sdr & (ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q )))

	.dataa(sdr),
	.datab(ram_rom_addr_reg_13),
	.datac(state_5),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h8000;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N26
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (sdr & (!ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q )))

	.dataa(sdr),
	.datab(ram_rom_addr_reg_13),
	.datac(state_5),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h2000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_mod_ram_rom (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg1,
	ram_rom_data_reg_0,
	ram_rom_addr_reg_13,
	ram_rom_addr_reg_0,
	ram_rom_addr_reg_1,
	ram_rom_addr_reg_2,
	ram_rom_addr_reg_3,
	ram_rom_addr_reg_4,
	ram_rom_addr_reg_5,
	ram_rom_addr_reg_6,
	ram_rom_addr_reg_7,
	ram_rom_addr_reg_8,
	ram_rom_addr_reg_9,
	ram_rom_addr_reg_10,
	ram_rom_addr_reg_11,
	ram_rom_addr_reg_12,
	ram_rom_data_reg_1,
	ram_rom_data_reg_2,
	ram_rom_data_reg_3,
	ram_rom_data_reg_4,
	ram_rom_data_reg_5,
	ram_rom_data_reg_6,
	ram_rom_data_reg_7,
	ram_rom_data_reg_8,
	ram_rom_data_reg_9,
	ram_rom_data_reg_10,
	ram_rom_data_reg_11,
	ram_rom_data_reg_12,
	ram_rom_data_reg_13,
	ram_rom_data_reg_14,
	ram_rom_data_reg_15,
	ram_rom_data_reg_16,
	ram_rom_data_reg_17,
	ram_rom_data_reg_18,
	ram_rom_data_reg_19,
	ram_rom_data_reg_20,
	ram_rom_data_reg_21,
	ram_rom_data_reg_22,
	ram_rom_data_reg_23,
	ram_rom_data_reg_24,
	ram_rom_data_reg_25,
	ram_rom_data_reg_26,
	ram_rom_data_reg_27,
	ram_rom_data_reg_28,
	ram_rom_data_reg_29,
	ram_rom_data_reg_30,
	ram_rom_data_reg_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	sdr,
	address_reg_b_0,
	altera_internal_jtag,
	state_4,
	ir_in,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_4_1,
	node_ena_1,
	clr,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	raw_tck,
	devpor,
	devclrn,
	devoe);
input 	ram_block3a32;
input 	ram_block3a0;
input 	ram_block3a33;
input 	ram_block3a1;
input 	ram_block3a34;
input 	ram_block3a2;
input 	ram_block3a35;
input 	ram_block3a3;
input 	ram_block3a36;
input 	ram_block3a4;
input 	ram_block3a37;
input 	ram_block3a5;
input 	ram_block3a38;
input 	ram_block3a6;
input 	ram_block3a39;
input 	ram_block3a7;
input 	ram_block3a40;
input 	ram_block3a8;
input 	ram_block3a41;
input 	ram_block3a9;
input 	ram_block3a42;
input 	ram_block3a10;
input 	ram_block3a43;
input 	ram_block3a11;
input 	ram_block3a44;
input 	ram_block3a12;
input 	ram_block3a45;
input 	ram_block3a13;
input 	ram_block3a46;
input 	ram_block3a14;
input 	ram_block3a47;
input 	ram_block3a15;
input 	ram_block3a48;
input 	ram_block3a16;
input 	ram_block3a49;
input 	ram_block3a17;
input 	ram_block3a50;
input 	ram_block3a18;
input 	ram_block3a51;
input 	ram_block3a19;
input 	ram_block3a52;
input 	ram_block3a20;
input 	ram_block3a53;
input 	ram_block3a21;
input 	ram_block3a54;
input 	ram_block3a22;
input 	ram_block3a55;
input 	ram_block3a23;
input 	ram_block3a56;
input 	ram_block3a24;
input 	ram_block3a57;
input 	ram_block3a25;
input 	ram_block3a58;
input 	ram_block3a26;
input 	ram_block3a59;
input 	ram_block3a27;
input 	ram_block3a60;
input 	ram_block3a28;
input 	ram_block3a61;
input 	ram_block3a29;
input 	ram_block3a62;
input 	ram_block3a30;
input 	ram_block3a63;
input 	ram_block3a31;
output 	is_in_use_reg1;
output 	ram_rom_data_reg_0;
output 	ram_rom_addr_reg_13;
output 	ram_rom_addr_reg_0;
output 	ram_rom_addr_reg_1;
output 	ram_rom_addr_reg_2;
output 	ram_rom_addr_reg_3;
output 	ram_rom_addr_reg_4;
output 	ram_rom_addr_reg_5;
output 	ram_rom_addr_reg_6;
output 	ram_rom_addr_reg_7;
output 	ram_rom_addr_reg_8;
output 	ram_rom_addr_reg_9;
output 	ram_rom_addr_reg_10;
output 	ram_rom_addr_reg_11;
output 	ram_rom_addr_reg_12;
output 	ram_rom_data_reg_1;
output 	ram_rom_data_reg_2;
output 	ram_rom_data_reg_3;
output 	ram_rom_data_reg_4;
output 	ram_rom_data_reg_5;
output 	ram_rom_data_reg_6;
output 	ram_rom_data_reg_7;
output 	ram_rom_data_reg_8;
output 	ram_rom_data_reg_9;
output 	ram_rom_data_reg_10;
output 	ram_rom_data_reg_11;
output 	ram_rom_data_reg_12;
output 	ram_rom_data_reg_13;
output 	ram_rom_data_reg_14;
output 	ram_rom_data_reg_15;
output 	ram_rom_data_reg_16;
output 	ram_rom_data_reg_17;
output 	ram_rom_data_reg_18;
output 	ram_rom_data_reg_19;
output 	ram_rom_data_reg_20;
output 	ram_rom_data_reg_21;
output 	ram_rom_data_reg_22;
output 	ram_rom_data_reg_23;
output 	ram_rom_data_reg_24;
output 	ram_rom_data_reg_25;
output 	ram_rom_data_reg_26;
output 	ram_rom_data_reg_27;
output 	ram_rom_data_reg_28;
output 	ram_rom_data_reg_29;
output 	ram_rom_data_reg_30;
output 	ram_rom_data_reg_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
output 	sdr;
input 	address_reg_b_0;
input 	altera_internal_jtag;
input 	state_4;
input 	[4:0] ir_in;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	raw_tck;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~9 ;
wire \Add1~10_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~10_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~12_combout ;
wire \is_in_use_reg~0_combout ;
wire \ram_rom_data_reg[0]~0_combout ;
wire \Add1~0_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~11_combout ;
wire \ram_rom_data_shift_cntr_reg[0]~6_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \ram_rom_data_shift_cntr_reg[1]~5_combout ;
wire \Add1~3 ;
wire \Add1~4_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~9_combout ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~7_combout ;
wire \Add1~6_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~8_combout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \process_0~2_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~4_combout ;
wire \ram_rom_data_reg[31]~32_combout ;
wire \ram_rom_addr_reg[0]~15 ;
wire \ram_rom_addr_reg[1]~17 ;
wire \ram_rom_addr_reg[2]~19 ;
wire \ram_rom_addr_reg[3]~21 ;
wire \ram_rom_addr_reg[4]~23 ;
wire \ram_rom_addr_reg[5]~25 ;
wire \ram_rom_addr_reg[6]~27 ;
wire \ram_rom_addr_reg[7]~29 ;
wire \ram_rom_addr_reg[8]~31 ;
wire \ram_rom_addr_reg[9]~33 ;
wire \ram_rom_addr_reg[10]~35 ;
wire \ram_rom_addr_reg[11]~37 ;
wire \ram_rom_addr_reg[12]~39 ;
wire \ram_rom_addr_reg[13]~40_combout ;
wire \process_0~3_combout ;
wire \ram_rom_addr_reg[5]~42_combout ;
wire \ram_rom_addr_reg[5]~43_combout ;
wire \ram_rom_addr_reg[0]~14_combout ;
wire \ram_rom_addr_reg[1]~16_combout ;
wire \ram_rom_addr_reg[2]~18_combout ;
wire \ram_rom_addr_reg[3]~20_combout ;
wire \ram_rom_addr_reg[4]~22_combout ;
wire \ram_rom_addr_reg[5]~24_combout ;
wire \ram_rom_addr_reg[6]~26_combout ;
wire \ram_rom_addr_reg[7]~28_combout ;
wire \ram_rom_addr_reg[8]~30_combout ;
wire \ram_rom_addr_reg[9]~32_combout ;
wire \ram_rom_addr_reg[10]~34_combout ;
wire \ram_rom_addr_reg[11]~36_combout ;
wire \ram_rom_addr_reg[12]~38_combout ;
wire \ram_rom_data_reg[1]~1_combout ;
wire \ram_rom_data_reg[2]~2_combout ;
wire \ram_rom_data_reg[3]~3_combout ;
wire \ram_rom_data_reg[4]~4_combout ;
wire \ram_rom_data_reg[5]~5_combout ;
wire \ram_rom_data_reg[6]~6_combout ;
wire \ram_rom_data_reg[7]~7_combout ;
wire \ram_rom_data_reg[8]~8_combout ;
wire \ram_rom_data_reg[9]~9_combout ;
wire \ram_rom_data_reg[10]~10_combout ;
wire \ram_rom_data_reg[11]~11_combout ;
wire \ram_rom_data_reg[12]~12_combout ;
wire \ram_rom_data_reg[13]~13_combout ;
wire \ram_rom_data_reg[14]~14_combout ;
wire \ram_rom_data_reg[15]~15_combout ;
wire \ram_rom_data_reg[16]~16_combout ;
wire \ram_rom_data_reg[17]~17_combout ;
wire \ram_rom_data_reg[18]~18_combout ;
wire \ram_rom_data_reg[19]~19_combout ;
wire \ram_rom_data_reg[20]~20_combout ;
wire \ram_rom_data_reg[21]~21_combout ;
wire \ram_rom_data_reg[22]~22_combout ;
wire \ram_rom_data_reg[23]~23_combout ;
wire \ram_rom_data_reg[24]~24_combout ;
wire \ram_rom_data_reg[25]~25_combout ;
wire \ram_rom_data_reg[26]~26_combout ;
wire \ram_rom_data_reg[27]~27_combout ;
wire \ram_rom_data_reg[28]~28_combout ;
wire \ram_rom_data_reg[29]~29_combout ;
wire \ram_rom_data_reg[30]~30_combout ;
wire \ram_rom_data_reg[31]~31_combout ;
wire \ir_loaded_address_reg[0]~feeder_combout ;
wire \process_0~0_combout ;
wire \process_0~1_combout ;
wire \ir_loaded_address_reg[1]~feeder_combout ;
wire \ir_loaded_address_reg[2]~feeder_combout ;
wire \ir_loaded_address_reg[3]~feeder_combout ;
wire \bypass_reg_out~0_combout ;
wire \bypass_reg_out~q ;
wire \tdo~0_combout ;
wire [5:0] ram_rom_data_shift_cntr_reg;
wire [3:0] \ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR ;


sld_rom_sr \ram_rom_logic_gen:name_gen:info_rom_sr (
	.WORD_SR_0(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.sdr(sdr),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.TCK(raw_tck),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X49_Y34_N20
cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N22
cycloneive_lcell_comb \Add1~10 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X49_Y34_N31
dffeas \ram_rom_data_shift_cntr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[5]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N30
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~10 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~10_combout ),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~10 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[5]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N10
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~12 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datab(ram_rom_data_shift_cntr_reg[0]),
	.datac(\Equal1~0_combout ),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~12 .lut_mask = 16'hD555;
defparam \ram_rom_data_shift_cntr_reg[5]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N21
dffeas is_in_use_reg(
	.clk(raw_tck),
	.d(\is_in_use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(ir_in[0]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(is_in_use_reg1),
	.prn(vcc));
// synopsys translate_off
defparam is_in_use_reg.is_wysiwyg = "true";
defparam is_in_use_reg.power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N25
dffeas \ram_rom_data_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[0]~0_combout ),
	.asdata(ram_rom_data_reg_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N29
dffeas \ram_rom_addr_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[13]~40_combout ),
	.asdata(altera_internal_jtag),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N3
dffeas \ram_rom_addr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[0]~14_combout ),
	.asdata(ram_rom_addr_reg_1),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N5
dffeas \ram_rom_addr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[1]~16_combout ),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N7
dffeas \ram_rom_addr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[2]~18_combout ),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N9
dffeas \ram_rom_addr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[3]~20_combout ),
	.asdata(ram_rom_addr_reg_4),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N11
dffeas \ram_rom_addr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[4]~22_combout ),
	.asdata(ram_rom_addr_reg_5),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N13
dffeas \ram_rom_addr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[5]~24_combout ),
	.asdata(ram_rom_addr_reg_6),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N15
dffeas \ram_rom_addr_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[6]~26_combout ),
	.asdata(ram_rom_addr_reg_7),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N17
dffeas \ram_rom_addr_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[7]~28_combout ),
	.asdata(ram_rom_addr_reg_8),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N19
dffeas \ram_rom_addr_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[8]~30_combout ),
	.asdata(ram_rom_addr_reg_9),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N21
dffeas \ram_rom_addr_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[9]~32_combout ),
	.asdata(ram_rom_addr_reg_10),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N23
dffeas \ram_rom_addr_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[10]~34_combout ),
	.asdata(ram_rom_addr_reg_11),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N25
dffeas \ram_rom_addr_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[11]~36_combout ),
	.asdata(ram_rom_addr_reg_12),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N27
dffeas \ram_rom_addr_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[12]~38_combout ),
	.asdata(ram_rom_addr_reg_13),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N23
dffeas \ram_rom_data_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[1]~1_combout ),
	.asdata(ram_rom_data_reg_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N13
dffeas \ram_rom_data_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[2]~2_combout ),
	.asdata(ram_rom_data_reg_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N15
dffeas \ram_rom_data_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[3]~3_combout ),
	.asdata(ram_rom_data_reg_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N9
dffeas \ram_rom_data_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[4]~4_combout ),
	.asdata(ram_rom_data_reg_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N11
dffeas \ram_rom_data_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[5]~5_combout ),
	.asdata(ram_rom_data_reg_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N29
dffeas \ram_rom_data_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[6]~6_combout ),
	.asdata(ram_rom_data_reg_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N31
dffeas \ram_rom_data_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[7]~7_combout ),
	.asdata(ram_rom_data_reg_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N5
dffeas \ram_rom_data_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[8]~8_combout ),
	.asdata(ram_rom_data_reg_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N27
dffeas \ram_rom_data_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[9]~9_combout ),
	.asdata(ram_rom_data_reg_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N1
dffeas \ram_rom_data_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[10]~10_combout ),
	.asdata(ram_rom_data_reg_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N5
dffeas \ram_rom_data_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[11]~11_combout ),
	.asdata(ram_rom_data_reg_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N17
dffeas \ram_rom_data_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[12]~12_combout ),
	.asdata(ram_rom_data_reg_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N31
dffeas \ram_rom_data_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[13]~13_combout ),
	.asdata(ram_rom_data_reg_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N25
dffeas \ram_rom_data_reg[14] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[14]~14_combout ),
	.asdata(ram_rom_data_reg_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_14),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[14] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N11
dffeas \ram_rom_data_reg[15] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[15]~15_combout ),
	.asdata(ram_rom_data_reg_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_15),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[15] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N13
dffeas \ram_rom_data_reg[16] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[16]~16_combout ),
	.asdata(ram_rom_data_reg_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_16),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[16] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N15
dffeas \ram_rom_data_reg[17] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[17]~17_combout ),
	.asdata(ram_rom_data_reg_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_17),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[17] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N9
dffeas \ram_rom_data_reg[18] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[18]~18_combout ),
	.asdata(ram_rom_data_reg_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_18),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[18] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N23
dffeas \ram_rom_data_reg[19] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[19]~19_combout ),
	.asdata(ram_rom_data_reg_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_19),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[19] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N29
dffeas \ram_rom_data_reg[20] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[20]~20_combout ),
	.asdata(ram_rom_data_reg_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_20),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[20] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N21
dffeas \ram_rom_data_reg[21] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[21]~21_combout ),
	.asdata(ram_rom_data_reg_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_21),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[21] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N1
dffeas \ram_rom_data_reg[22] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[22]~22_combout ),
	.asdata(ram_rom_data_reg_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_22),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[22] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N19
dffeas \ram_rom_data_reg[23] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[23]~23_combout ),
	.asdata(ram_rom_data_reg_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_23),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[23] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N27
dffeas \ram_rom_data_reg[24] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[24]~24_combout ),
	.asdata(ram_rom_data_reg_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_24),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[24] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N17
dffeas \ram_rom_data_reg[25] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[25]~25_combout ),
	.asdata(ram_rom_data_reg_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_25),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[25] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N15
dffeas \ram_rom_data_reg[26] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[26]~26_combout ),
	.asdata(ram_rom_data_reg_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_26),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[26] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N29
dffeas \ram_rom_data_reg[27] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[27]~27_combout ),
	.asdata(ram_rom_data_reg_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_27),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[27] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N11
dffeas \ram_rom_data_reg[28] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[28]~28_combout ),
	.asdata(ram_rom_data_reg_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_28),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[28] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N9
dffeas \ram_rom_data_reg[29] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[29]~29_combout ),
	.asdata(ram_rom_data_reg_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_29),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[29] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N23
dffeas \ram_rom_data_reg[30] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[30]~30_combout ),
	.asdata(ram_rom_data_reg_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_30),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[30] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N13
dffeas \ram_rom_data_reg[31] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[31]~31_combout ),
	.asdata(altera_internal_jtag),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_31),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[31] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N9
dffeas \ir_loaded_address_reg[0] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[0] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N11
dffeas \ir_loaded_address_reg[1] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[1] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N5
dffeas \ir_loaded_address_reg[2] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[2] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N23
dffeas \ir_loaded_address_reg[3] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[3] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N0
cycloneive_lcell_comb \tdo~1 (
	.dataa(\tdo~0_combout ),
	.datab(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.datac(ir_in[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(tdo),
	.cout());
// synopsys translate_off
defparam \tdo~1 .lut_mask = 16'hCACA;
defparam \tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N10
cycloneive_lcell_comb \sdr~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(node_ena_1),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(sdr),
	.cout());
// synopsys translate_off
defparam \sdr~0 .lut_mask = 16'h00F0;
defparam \sdr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N20
cycloneive_lcell_comb \is_in_use_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(is_in_use_reg1),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\is_in_use_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \is_in_use_reg~0 .lut_mask = 16'h00F0;
defparam \is_in_use_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N24
cycloneive_lcell_comb \ram_rom_data_reg[0]~0 (
	.dataa(ram_block3a32),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~0 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N12
cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h33CC;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N28
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~11 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datab(ram_rom_data_shift_cntr_reg[0]),
	.datac(\Equal1~0_combout ),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~11 .lut_mask = 16'h1555;
defparam \ram_rom_data_shift_cntr_reg[5]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N2
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[0]~6 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0]~6 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N3
dffeas \ram_rom_data_shift_cntr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N14
cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h3C3F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N0
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[1]~5 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datab(\Add1~2_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1]~5 .lut_mask = 16'h08D8;
defparam \ram_rom_data_shift_cntr_reg[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N1
dffeas \ram_rom_data_shift_cntr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N16
cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hC30C;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N8
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~9 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~4_combout ),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~9 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N9
dffeas \ram_rom_data_shift_cntr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N18
cycloneive_lcell_comb \Add1~6 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N24
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~7 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~8_combout ),
	.datac(ram_rom_data_shift_cntr_reg[4]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~7 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N25
dffeas \ram_rom_data_shift_cntr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[4]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N6
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~8 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~6_combout ),
	.datac(ram_rom_data_shift_cntr_reg[3]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~8 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N7
dffeas \ram_rom_data_shift_cntr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N4
cycloneive_lcell_comb \Equal1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(ram_rom_data_shift_cntr_reg[3]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h4000;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N26
cycloneive_lcell_comb \Equal1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\Equal1~0_combout ),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'hF000;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N26
cycloneive_lcell_comb \process_0~2 (
	.dataa(\Equal1~1_combout ),
	.datab(ir_in[3]),
	.datac(irf_reg_1_1),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~2 .lut_mask = 16'h1333;
defparam \process_0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N14
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~4 (
	.dataa(irf_reg_1_1),
	.datab(sdr),
	.datac(state_4),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~4 .lut_mask = 16'hC080;
defparam \ram_rom_data_shift_cntr_reg[5]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N18
cycloneive_lcell_comb \ram_rom_data_reg[31]~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\process_0~2_combout ),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~32_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~32 .lut_mask = 16'hFF0F;
defparam \ram_rom_data_reg[31]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N2
cycloneive_lcell_comb \ram_rom_addr_reg[0]~14 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[0]~14_combout ),
	.cout(\ram_rom_addr_reg[0]~15 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[0]~14 .lut_mask = 16'h33CC;
defparam \ram_rom_addr_reg[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N4
cycloneive_lcell_comb \ram_rom_addr_reg[1]~16 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[0]~15 ),
	.combout(\ram_rom_addr_reg[1]~16_combout ),
	.cout(\ram_rom_addr_reg[1]~17 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~16 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[1]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N6
cycloneive_lcell_comb \ram_rom_addr_reg[2]~18 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[1]~17 ),
	.combout(\ram_rom_addr_reg[2]~18_combout ),
	.cout(\ram_rom_addr_reg[2]~19 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~18 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[2]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N8
cycloneive_lcell_comb \ram_rom_addr_reg[3]~20 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[2]~19 ),
	.combout(\ram_rom_addr_reg[3]~20_combout ),
	.cout(\ram_rom_addr_reg[3]~21 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[3]~20 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[3]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N10
cycloneive_lcell_comb \ram_rom_addr_reg[4]~22 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[3]~21 ),
	.combout(\ram_rom_addr_reg[4]~22_combout ),
	.cout(\ram_rom_addr_reg[4]~23 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~22 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[4]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N12
cycloneive_lcell_comb \ram_rom_addr_reg[5]~24 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[4]~23 ),
	.combout(\ram_rom_addr_reg[5]~24_combout ),
	.cout(\ram_rom_addr_reg[5]~25 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~24 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[5]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N14
cycloneive_lcell_comb \ram_rom_addr_reg[6]~26 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[5]~25 ),
	.combout(\ram_rom_addr_reg[6]~26_combout ),
	.cout(\ram_rom_addr_reg[6]~27 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~26 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[6]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N16
cycloneive_lcell_comb \ram_rom_addr_reg[7]~28 (
	.dataa(ram_rom_addr_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[6]~27 ),
	.combout(\ram_rom_addr_reg[7]~28_combout ),
	.cout(\ram_rom_addr_reg[7]~29 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~28 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[7]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N18
cycloneive_lcell_comb \ram_rom_addr_reg[8]~30 (
	.dataa(ram_rom_addr_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[7]~29 ),
	.combout(\ram_rom_addr_reg[8]~30_combout ),
	.cout(\ram_rom_addr_reg[8]~31 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[8]~30 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[8]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N20
cycloneive_lcell_comb \ram_rom_addr_reg[9]~32 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[8]~31 ),
	.combout(\ram_rom_addr_reg[9]~32_combout ),
	.cout(\ram_rom_addr_reg[9]~33 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~32 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[9]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N22
cycloneive_lcell_comb \ram_rom_addr_reg[10]~34 (
	.dataa(ram_rom_addr_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[9]~33 ),
	.combout(\ram_rom_addr_reg[10]~34_combout ),
	.cout(\ram_rom_addr_reg[10]~35 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[10]~34 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[10]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N24
cycloneive_lcell_comb \ram_rom_addr_reg[11]~36 (
	.dataa(ram_rom_addr_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[10]~35 ),
	.combout(\ram_rom_addr_reg[11]~36_combout ),
	.cout(\ram_rom_addr_reg[11]~37 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[11]~36 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[11]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N26
cycloneive_lcell_comb \ram_rom_addr_reg[12]~38 (
	.dataa(ram_rom_addr_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[11]~37 ),
	.combout(\ram_rom_addr_reg[12]~38_combout ),
	.cout(\ram_rom_addr_reg[12]~39 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[12]~38 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[12]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N28
cycloneive_lcell_comb \ram_rom_addr_reg[13]~40 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_13),
	.datac(gnd),
	.datad(gnd),
	.cin(\ram_rom_addr_reg[12]~39 ),
	.combout(\ram_rom_addr_reg[13]~40_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[13]~40 .lut_mask = 16'h3C3C;
defparam \ram_rom_addr_reg[13]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N28
cycloneive_lcell_comb \process_0~3 (
	.dataa(ir_in[3]),
	.datab(node_ena_1),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\process_0~3_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~3 .lut_mask = 16'h0080;
defparam \process_0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N30
cycloneive_lcell_comb \ram_rom_addr_reg[5]~42 (
	.dataa(\process_0~3_combout ),
	.datab(irf_reg_1_1),
	.datac(\Equal1~1_combout ),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[5]~42_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~42 .lut_mask = 16'hAAEA;
defparam \ram_rom_addr_reg[5]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N0
cycloneive_lcell_comb \ram_rom_addr_reg[5]~43 (
	.dataa(\ram_rom_addr_reg[5]~42_combout ),
	.datab(sdr),
	.datac(state_8),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[5]~43_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~43 .lut_mask = 16'hEAAA;
defparam \ram_rom_addr_reg[5]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N22
cycloneive_lcell_comb \ram_rom_data_reg[1]~1 (
	.dataa(ram_block3a33),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_rom_data_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[1]~1 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N12
cycloneive_lcell_comb \ram_rom_data_reg[2]~2 (
	.dataa(ram_block3a34),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a2),
	.cin(gnd),
	.combout(\ram_rom_data_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[2]~2 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N14
cycloneive_lcell_comb \ram_rom_data_reg[3]~3 (
	.dataa(ram_block3a35),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a3),
	.cin(gnd),
	.combout(\ram_rom_data_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[3]~3 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N8
cycloneive_lcell_comb \ram_rom_data_reg[4]~4 (
	.dataa(ram_block3a4),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a36),
	.cin(gnd),
	.combout(\ram_rom_data_reg[4]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[4]~4 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N10
cycloneive_lcell_comb \ram_rom_data_reg[5]~5 (
	.dataa(ram_block3a5),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a37),
	.cin(gnd),
	.combout(\ram_rom_data_reg[5]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[5]~5 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N28
cycloneive_lcell_comb \ram_rom_data_reg[6]~6 (
	.dataa(ram_block3a6),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a38),
	.cin(gnd),
	.combout(\ram_rom_data_reg[6]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[6]~6 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N30
cycloneive_lcell_comb \ram_rom_data_reg[7]~7 (
	.dataa(ram_block3a39),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a7),
	.cin(gnd),
	.combout(\ram_rom_data_reg[7]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[7]~7 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N4
cycloneive_lcell_comb \ram_rom_data_reg[8]~8 (
	.dataa(ram_block3a8),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a40),
	.cin(gnd),
	.combout(\ram_rom_data_reg[8]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[8]~8 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N26
cycloneive_lcell_comb \ram_rom_data_reg[9]~9 (
	.dataa(ram_block3a41),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a9),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~9 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N0
cycloneive_lcell_comb \ram_rom_data_reg[10]~10 (
	.dataa(ram_block3a10),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a42),
	.cin(gnd),
	.combout(\ram_rom_data_reg[10]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[10]~10 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N4
cycloneive_lcell_comb \ram_rom_data_reg[11]~11 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a43),
	.datac(gnd),
	.datad(ram_block3a11),
	.cin(gnd),
	.combout(\ram_rom_data_reg[11]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[11]~11 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N16
cycloneive_lcell_comb \ram_rom_data_reg[12]~12 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a44),
	.datac(gnd),
	.datad(ram_block3a12),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~12 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N30
cycloneive_lcell_comb \ram_rom_data_reg[13]~13 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a45),
	.datac(gnd),
	.datad(ram_block3a13),
	.cin(gnd),
	.combout(\ram_rom_data_reg[13]~13_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[13]~13 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N24
cycloneive_lcell_comb \ram_rom_data_reg[14]~14 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a14),
	.datac(gnd),
	.datad(ram_block3a46),
	.cin(gnd),
	.combout(\ram_rom_data_reg[14]~14_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[14]~14 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N10
cycloneive_lcell_comb \ram_rom_data_reg[15]~15 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a47),
	.datac(gnd),
	.datad(ram_block3a15),
	.cin(gnd),
	.combout(\ram_rom_data_reg[15]~15_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[15]~15 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N12
cycloneive_lcell_comb \ram_rom_data_reg[16]~16 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a48),
	.datac(gnd),
	.datad(ram_block3a16),
	.cin(gnd),
	.combout(\ram_rom_data_reg[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[16]~16 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N14
cycloneive_lcell_comb \ram_rom_data_reg[17]~17 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a17),
	.datac(gnd),
	.datad(ram_block3a49),
	.cin(gnd),
	.combout(\ram_rom_data_reg[17]~17_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[17]~17 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N8
cycloneive_lcell_comb \ram_rom_data_reg[18]~18 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a18),
	.datac(gnd),
	.datad(ram_block3a50),
	.cin(gnd),
	.combout(\ram_rom_data_reg[18]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[18]~18 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N22
cycloneive_lcell_comb \ram_rom_data_reg[19]~19 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a51),
	.datac(gnd),
	.datad(ram_block3a19),
	.cin(gnd),
	.combout(\ram_rom_data_reg[19]~19_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[19]~19 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N28
cycloneive_lcell_comb \ram_rom_data_reg[20]~20 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a20),
	.datac(gnd),
	.datad(ram_block3a52),
	.cin(gnd),
	.combout(\ram_rom_data_reg[20]~20_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[20]~20 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N20
cycloneive_lcell_comb \ram_rom_data_reg[21]~21 (
	.dataa(ram_block3a21),
	.datab(ram_block3a53),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~21 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N0
cycloneive_lcell_comb \ram_rom_data_reg[22]~22 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a22),
	.datac(gnd),
	.datad(ram_block3a54),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~22_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~22 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N18
cycloneive_lcell_comb \ram_rom_data_reg[23]~23 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a23),
	.datac(gnd),
	.datad(ram_block3a55),
	.cin(gnd),
	.combout(\ram_rom_data_reg[23]~23_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[23]~23 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N26
cycloneive_lcell_comb \ram_rom_data_reg[24]~24 (
	.dataa(ram_block3a24),
	.datab(ram_block3a56),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[24]~24_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[24]~24 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N16
cycloneive_lcell_comb \ram_rom_data_reg[25]~25 (
	.dataa(ram_block3a25),
	.datab(ram_block3a57),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[25]~25_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[25]~25 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N14
cycloneive_lcell_comb \ram_rom_data_reg[26]~26 (
	.dataa(ram_block3a26),
	.datab(ram_block3a58),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~26_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~26 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N28
cycloneive_lcell_comb \ram_rom_data_reg[27]~27 (
	.dataa(ram_block3a59),
	.datab(ram_block3a27),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[27]~27_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[27]~27 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N10
cycloneive_lcell_comb \ram_rom_data_reg[28]~28 (
	.dataa(ram_block3a60),
	.datab(ram_block3a28),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[28]~28_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[28]~28 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N8
cycloneive_lcell_comb \ram_rom_data_reg[29]~29 (
	.dataa(ram_block3a29),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a61),
	.cin(gnd),
	.combout(\ram_rom_data_reg[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[29]~29 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N22
cycloneive_lcell_comb \ram_rom_data_reg[30]~30 (
	.dataa(ram_block3a62),
	.datab(ram_block3a30),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[30]~30 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N12
cycloneive_lcell_comb \ram_rom_data_reg[31]~31 (
	.dataa(ram_block3a63),
	.datab(ram_block3a31),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~31_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~31 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N8
cycloneive_lcell_comb \ir_loaded_address_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_0),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N14
cycloneive_lcell_comb \process_0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ir_in[0]),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~0 .lut_mask = 16'hFFF0;
defparam \process_0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N12
cycloneive_lcell_comb \process_0~1 (
	.dataa(ir_in[3]),
	.datab(node_ena_1),
	.datac(state_5),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~1 .lut_mask = 16'h0080;
defparam \process_0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N10
cycloneive_lcell_comb \ir_loaded_address_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_1),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N4
cycloneive_lcell_comb \ir_loaded_address_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_2),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N22
cycloneive_lcell_comb \ir_loaded_address_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_3),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N0
cycloneive_lcell_comb \bypass_reg_out~0 (
	.dataa(altera_internal_jtag),
	.datab(gnd),
	.datac(\bypass_reg_out~q ),
	.datad(node_ena_1),
	.cin(gnd),
	.combout(\bypass_reg_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \bypass_reg_out~0 .lut_mask = 16'hAAF0;
defparam \bypass_reg_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y37_N1
dffeas bypass_reg_out(
	.clk(raw_tck),
	.d(\bypass_reg_out~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bypass_reg_out~q ),
	.prn(vcc));
// synopsys translate_off
defparam bypass_reg_out.is_wysiwyg = "true";
defparam bypass_reg_out.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N30
cycloneive_lcell_comb \tdo~0 (
	.dataa(irf_reg_1_1),
	.datab(ram_rom_data_reg_0),
	.datac(\bypass_reg_out~q ),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \tdo~0 .lut_mask = 16'hCCD8;
defparam \tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_rom_sr (
	WORD_SR_0,
	sdr,
	altera_internal_jtag,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	TCK,
	devpor,
	devclrn,
	devoe);
output 	WORD_SR_0;
input 	sdr;
input 	altera_internal_jtag;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	TCK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \word_counter[3]~15_combout ;
wire \WORD_SR~7_combout ;
wire \WORD_SR~8_combout ;
wire \WORD_SR~10_combout ;
wire \WORD_SR~13_combout ;
wire \WORD_SR~14_combout ;
wire \WORD_SR~15_combout ;
wire \clear_signal~combout ;
wire \word_counter[0]~7_combout ;
wire \word_counter[1]~9_combout ;
wire \word_counter[1]~14_combout ;
wire \word_counter[1]~13_combout ;
wire \word_counter[1]~19_combout ;
wire \word_counter[0]~8 ;
wire \word_counter[1]~10 ;
wire \word_counter[2]~11_combout ;
wire \word_counter[2]~12 ;
wire \word_counter[3]~16 ;
wire \word_counter[4]~17_combout ;
wire \WORD_SR~2_combout ;
wire \WORD_SR~11_combout ;
wire \WORD_SR~12_combout ;
wire \WORD_SR[2]~6_combout ;
wire \WORD_SR~9_combout ;
wire \WORD_SR~3_combout ;
wire \WORD_SR~4_combout ;
wire \WORD_SR~5_combout ;
wire [4:0] word_counter;
wire [3:0] WORD_SR;


// Location: FF_X47_Y37_N11
dffeas \word_counter[3] (
	.clk(TCK),
	.d(\word_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[3]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[3] .is_wysiwyg = "true";
defparam \word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N10
cycloneive_lcell_comb \word_counter[3]~15 (
	.dataa(word_counter[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[2]~12 ),
	.combout(\word_counter[3]~15_combout ),
	.cout(\word_counter[3]~16 ));
// synopsys translate_off
defparam \word_counter[3]~15 .lut_mask = 16'h5A5F;
defparam \word_counter[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N16
cycloneive_lcell_comb \WORD_SR~7 (
	.dataa(word_counter[1]),
	.datab(state_4),
	.datac(word_counter[0]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~7 .lut_mask = 16'h0203;
defparam \WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N26
cycloneive_lcell_comb \WORD_SR~8 (
	.dataa(gnd),
	.datab(\WORD_SR~7_combout ),
	.datac(word_counter[2]),
	.datad(word_counter[3]),
	.cin(gnd),
	.combout(\WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~8 .lut_mask = 16'h000C;
defparam \WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N23
dffeas \WORD_SR[3] (
	.clk(TCK),
	.d(\WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[3]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[3] .is_wysiwyg = "true";
defparam \WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N30
cycloneive_lcell_comb \WORD_SR~10 (
	.dataa(word_counter[1]),
	.datab(word_counter[2]),
	.datac(word_counter[0]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~10 .lut_mask = 16'hF784;
defparam \WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N18
cycloneive_lcell_comb \WORD_SR~13 (
	.dataa(word_counter[3]),
	.datab(word_counter[4]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~13 .lut_mask = 16'h2000;
defparam \WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N20
cycloneive_lcell_comb \WORD_SR~14 (
	.dataa(altera_internal_jtag),
	.datab(state_4),
	.datac(word_counter[0]),
	.datad(\WORD_SR~13_combout ),
	.cin(gnd),
	.combout(\WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~14 .lut_mask = 16'h8B88;
defparam \WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N22
cycloneive_lcell_comb \WORD_SR~15 (
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(state_8),
	.datad(\WORD_SR~14_combout ),
	.cin(gnd),
	.combout(\WORD_SR~15_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~15 .lut_mask = 16'h5F00;
defparam \WORD_SR~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N21
dffeas \WORD_SR[0] (
	.clk(TCK),
	.d(\WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR_0),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[0] .is_wysiwyg = "true";
defparam \WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N16
cycloneive_lcell_comb clear_signal(
	.dataa(gnd),
	.datab(gnd),
	.datac(state_8),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam clear_signal.lut_mask = 16'hF000;
defparam clear_signal.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N4
cycloneive_lcell_comb \word_counter[0]~7 (
	.dataa(gnd),
	.datab(word_counter[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\word_counter[0]~7_combout ),
	.cout(\word_counter[0]~8 ));
// synopsys translate_off
defparam \word_counter[0]~7 .lut_mask = 16'h33CC;
defparam \word_counter[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N6
cycloneive_lcell_comb \word_counter[1]~9 (
	.dataa(word_counter[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[0]~8 ),
	.combout(\word_counter[1]~9_combout ),
	.cout(\word_counter[1]~10 ));
// synopsys translate_off
defparam \word_counter[1]~9 .lut_mask = 16'h5A5F;
defparam \word_counter[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N8
cycloneive_lcell_comb \word_counter[1]~14 (
	.dataa(sdr),
	.datab(state_3),
	.datac(state_4),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\word_counter[1]~14_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[1]~14 .lut_mask = 16'hFF08;
defparam \word_counter[1]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y37_N7
dffeas \word_counter[1] (
	.clk(TCK),
	.d(\word_counter[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[1]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[1] .is_wysiwyg = "true";
defparam \word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N28
cycloneive_lcell_comb \word_counter[1]~13 (
	.dataa(word_counter[3]),
	.datab(word_counter[4]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\word_counter[1]~13_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[1]~13 .lut_mask = 16'hFFBF;
defparam \word_counter[1]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N2
cycloneive_lcell_comb \word_counter[1]~19 (
	.dataa(state_8),
	.datab(virtual_ir_scan_reg),
	.datac(word_counter[0]),
	.datad(\word_counter[1]~13_combout ),
	.cin(gnd),
	.combout(\word_counter[1]~19_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[1]~19 .lut_mask = 16'h888F;
defparam \word_counter[1]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y37_N5
dffeas \word_counter[0] (
	.clk(TCK),
	.d(\word_counter[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[0]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[0] .is_wysiwyg = "true";
defparam \word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N8
cycloneive_lcell_comb \word_counter[2]~11 (
	.dataa(gnd),
	.datab(word_counter[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[1]~10 ),
	.combout(\word_counter[2]~11_combout ),
	.cout(\word_counter[2]~12 ));
// synopsys translate_off
defparam \word_counter[2]~11 .lut_mask = 16'hC30C;
defparam \word_counter[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X47_Y37_N9
dffeas \word_counter[2] (
	.clk(TCK),
	.d(\word_counter[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[2]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[2] .is_wysiwyg = "true";
defparam \word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N12
cycloneive_lcell_comb \word_counter[4]~17 (
	.dataa(word_counter[4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\word_counter[3]~16 ),
	.combout(\word_counter[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~17 .lut_mask = 16'hA5A5;
defparam \word_counter[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X47_Y37_N13
dffeas \word_counter[4] (
	.clk(TCK),
	.d(\word_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[4]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[4] .is_wysiwyg = "true";
defparam \word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N14
cycloneive_lcell_comb \WORD_SR~2 (
	.dataa(word_counter[3]),
	.datab(word_counter[4]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~2_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~2 .lut_mask = 16'h2025;
defparam \WORD_SR~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N24
cycloneive_lcell_comb \WORD_SR~11 (
	.dataa(\WORD_SR~10_combout ),
	.datab(\WORD_SR~2_combout ),
	.datac(word_counter[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~11 .lut_mask = 16'hA4A4;
defparam \WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N18
cycloneive_lcell_comb \WORD_SR~12 (
	.dataa(WORD_SR[3]),
	.datab(\WORD_SR~11_combout ),
	.datac(state_4),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~12 .lut_mask = 16'h00AC;
defparam \WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N4
cycloneive_lcell_comb \WORD_SR[2]~6 (
	.dataa(sdr),
	.datab(state_3),
	.datac(state_4),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR[2]~6_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR[2]~6 .lut_mask = 16'hFFA8;
defparam \WORD_SR[2]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N19
dffeas \WORD_SR[2] (
	.clk(TCK),
	.d(\WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[2]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[2] .is_wysiwyg = "true";
defparam \WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N6
cycloneive_lcell_comb \WORD_SR~9 (
	.dataa(\WORD_SR~8_combout ),
	.datab(\clear_signal~combout ),
	.datac(state_4),
	.datad(WORD_SR[2]),
	.cin(gnd),
	.combout(\WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~9 .lut_mask = 16'h3222;
defparam \WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N7
dffeas \WORD_SR[1] (
	.clk(TCK),
	.d(\WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[1]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[1] .is_wysiwyg = "true";
defparam \WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N22
cycloneive_lcell_comb \WORD_SR~3 (
	.dataa(word_counter[1]),
	.datab(word_counter[2]),
	.datac(word_counter[0]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~3_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~3 .lut_mask = 16'hAB08;
defparam \WORD_SR~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N2
cycloneive_lcell_comb \WORD_SR~4 (
	.dataa(gnd),
	.datab(\WORD_SR~3_combout ),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~4_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~4 .lut_mask = 16'hCCC0;
defparam \WORD_SR~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N20
cycloneive_lcell_comb \WORD_SR~5 (
	.dataa(WORD_SR[1]),
	.datab(\clear_signal~combout ),
	.datac(state_4),
	.datad(\WORD_SR~4_combout ),
	.cin(gnd),
	.combout(\WORD_SR~5_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~5 .lut_mask = 16'h2320;
defparam \WORD_SR~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module singlecycle (
	PC_29,
	PC_28,
	PC_31,
	PC_30,
	dpifhalt,
	ramiframload_0,
	LessThan1,
	PC_1,
	daddr_1,
	ruifdWEN_r,
	ruifdREN_r,
	daddr_0,
	PC_0,
	daddr_3,
	PC_3,
	daddr_2,
	PC_2,
	daddr_5,
	PC_5,
	daddr_4,
	PC_4,
	daddr_7,
	PC_7,
	daddr_6,
	PC_6,
	always0,
	daddr_9,
	PC_9,
	PC_8,
	daddr_8,
	daddr_11,
	PC_11,
	daddr_10,
	PC_10,
	daddr_13,
	PC_13,
	daddr_12,
	PC_12,
	daddr_15,
	PC_15,
	daddr_14,
	PC_14,
	always01,
	PC_17,
	daddr_17,
	daddr_16,
	PC_16,
	daddr_19,
	PC_19,
	daddr_18,
	PC_18,
	PC_21,
	daddr_21,
	PC_20,
	daddr_20,
	daddr_23,
	PC_23,
	daddr_22,
	PC_22,
	daddr_25,
	PC_25,
	daddr_24,
	PC_24,
	daddr_27,
	PC_27,
	daddr_26,
	PC_26,
	daddr_29,
	daddr_28,
	daddr_31,
	daddr_30,
	always02,
	always03,
	ramiframload_01,
	always1,
	ramiframload_1,
	ramiframload_2,
	ramiframload_21,
	ramiframload_3,
	ramiframload_4,
	ramiframload_41,
	ramiframload_5,
	ramiframload_51,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_161,
	ramiframload_17,
	ramiframload_171,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_211,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_261,
	ramiframload_27,
	ramiframload_271,
	ramiframload_28,
	ramiframload_281,
	ramiframload_29,
	ramiframload_291,
	ramiframload_30,
	ramiframload_301,
	ramiframload_31,
	ramiframload_311,
	Mux63,
	Mux631,
	dcifimemload_20,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux36,
	Mux361,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux44,
	Mux441,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	Mux49,
	Mux491,
	Mux50,
	Mux501,
	Mux51,
	Mux511,
	Mux52,
	Mux521,
	Mux53,
	Mux531,
	Mux54,
	Mux541,
	Mux55,
	Mux551,
	Mux56,
	Mux561,
	Mux57,
	Mux571,
	Mux58,
	Mux581,
	Mux59,
	Mux591,
	Mux60,
	Mux601,
	Mux61,
	Mux611,
	Mux62,
	Mux621,
	Mux32,
	Mux321,
	nRST,
	CLK,
	nRST1,
	dpifhalt1,
	devpor,
	devclrn,
	devoe);
output 	PC_29;
output 	PC_28;
output 	PC_31;
output 	PC_30;
output 	dpifhalt;
input 	ramiframload_0;
input 	LessThan1;
output 	PC_1;
output 	daddr_1;
output 	ruifdWEN_r;
output 	ruifdREN_r;
output 	daddr_0;
output 	PC_0;
output 	daddr_3;
output 	PC_3;
output 	daddr_2;
output 	PC_2;
output 	daddr_5;
output 	PC_5;
output 	daddr_4;
output 	PC_4;
output 	daddr_7;
output 	PC_7;
output 	daddr_6;
output 	PC_6;
input 	always0;
output 	daddr_9;
output 	PC_9;
output 	PC_8;
output 	daddr_8;
output 	daddr_11;
output 	PC_11;
output 	daddr_10;
output 	PC_10;
output 	daddr_13;
output 	PC_13;
output 	daddr_12;
output 	PC_12;
output 	daddr_15;
output 	PC_15;
output 	daddr_14;
output 	PC_14;
input 	always01;
output 	PC_17;
output 	daddr_17;
output 	daddr_16;
output 	PC_16;
output 	daddr_19;
output 	PC_19;
output 	daddr_18;
output 	PC_18;
output 	PC_21;
output 	daddr_21;
output 	PC_20;
output 	daddr_20;
output 	daddr_23;
output 	PC_23;
output 	daddr_22;
output 	PC_22;
output 	daddr_25;
output 	PC_25;
output 	daddr_24;
output 	PC_24;
output 	daddr_27;
output 	PC_27;
output 	daddr_26;
output 	PC_26;
output 	daddr_29;
output 	daddr_28;
output 	daddr_31;
output 	daddr_30;
input 	always02;
input 	always03;
input 	ramiframload_01;
input 	always1;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_21;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_41;
input 	ramiframload_5;
input 	ramiframload_51;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_161;
input 	ramiframload_17;
input 	ramiframload_171;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_211;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_261;
input 	ramiframload_27;
input 	ramiframload_271;
input 	ramiframload_28;
input 	ramiframload_281;
input 	ramiframload_29;
input 	ramiframload_291;
input 	ramiframload_30;
input 	ramiframload_301;
input 	ramiframload_31;
input 	ramiframload_311;
output 	Mux63;
output 	Mux631;
output 	dcifimemload_20;
output 	Mux33;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux36;
output 	Mux361;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux41;
output 	Mux411;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux44;
output 	Mux441;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux48;
output 	Mux481;
output 	Mux49;
output 	Mux491;
output 	Mux50;
output 	Mux501;
output 	Mux51;
output 	Mux511;
output 	Mux52;
output 	Mux521;
output 	Mux53;
output 	Mux531;
output 	Mux54;
output 	Mux541;
output 	Mux55;
output 	Mux551;
output 	Mux56;
output 	Mux561;
output 	Mux57;
output 	Mux571;
output 	Mux58;
output 	Mux581;
output 	Mux59;
output 	Mux591;
output 	Mux60;
output 	Mux601;
output 	Mux61;
output 	Mux611;
output 	Mux62;
output 	Mux621;
output 	Mux32;
output 	Mux321;
input 	nRST;
input 	CLK;
input 	nRST1;
output 	dpifhalt1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \CC|ccif.iwait[0]~0_combout ;
wire \CM|dcif.imemload[26]~0_combout ;
wire \CM|dcif.imemload[27]~1_combout ;
wire \CM|dcif.imemload[28]~2_combout ;
wire \CM|dcif.imemload[29]~3_combout ;
wire \CM|dcif.imemload[30]~4_combout ;
wire \CM|dcif.imemload[31]~5_combout ;
wire \CM|dcif.ihit~0_combout ;
wire \CM|dcif.imemload[19]~6_combout ;
wire \CM|dcif.imemload[18]~7_combout ;
wire \CM|dcif.imemload[16]~8_combout ;
wire \CM|dcif.imemload[17]~9_combout ;
wire \CM|dcif.imemload[24]~11_combout ;
wire \CM|dcif.imemload[23]~12_combout ;
wire \CM|dcif.imemload[21]~13_combout ;
wire \CM|dcif.imemload[22]~14_combout ;
wire \CM|dcif.imemload[25]~15_combout ;
wire \CM|dcif.imemload[3]~16_combout ;
wire \CM|dcif.imemload[4]~17_combout ;
wire \CM|dcif.imemload[2]~18_combout ;
wire \CM|dcif.imemload[5]~19_combout ;
wire \CM|dcif.imemload[0]~20_combout ;
wire \CM|dcif.imemload[1]~21_combout ;
wire \CM|dcif.imemload[15]~22_combout ;
wire \CM|dcif.imemload[14]~23_combout ;
wire \CM|dcif.imemload[13]~24_combout ;
wire \CM|dcif.imemload[12]~25_combout ;
wire \CM|dcif.imemload[11]~26_combout ;
wire \CM|dcif.imemload[10]~27_combout ;
wire \CM|dcif.imemload[9]~28_combout ;
wire \CM|dcif.imemload[8]~29_combout ;
wire \CM|dcif.imemload[7]~30_combout ;
wire \CM|dcif.imemload[6]~31_combout ;
wire \DP|cu|Selector0~2_combout ;
wire \DP|ALU|Mux1~7_combout ;
wire \DP|ALU|Mux31~0_combout ;
wire \DP|ALU|Mux1~8_combout ;
wire \DP|ALU|Mux0~13_combout ;
wire \DP|ALU|Mux0~14_combout ;
wire \DP|ALU|Mux24~9_combout ;
wire \DP|ALU|Mux25~5_combout ;
wire \DP|ALU|Mux26~5_combout ;
wire \DP|ALU|Mux27~5_combout ;
wire \DP|ALU|Mux4~6_combout ;
wire \DP|ALU|Mux5~6_combout ;
wire \DP|ALU|Mux6~16_combout ;
wire \DP|ALU|Mux7~6_combout ;
wire \DP|ALU|Mux3~7_combout ;
wire \DP|ALU|Mux2~11_combout ;
wire \DP|ALU|Mux23~7_combout ;
wire \DP|ALU|Mux23~8_combout ;
wire \DP|ALU|Mux22~5_combout ;
wire \DP|ALU|Mux22~6_combout ;
wire \DP|ALU|Mux21~5_combout ;
wire \DP|ALU|Mux21~6_combout ;
wire \DP|ALU|Mux20~5_combout ;
wire \DP|ALU|Mux20~6_combout ;
wire \DP|ALU|Mux19~5_combout ;
wire \DP|ALU|Mux19~6_combout ;
wire \DP|ALU|Mux18~8_combout ;
wire \DP|ALU|Mux18~9_combout ;
wire \DP|ALU|Mux17~5_combout ;
wire \DP|ALU|Mux17~6_combout ;
wire \DP|ALU|Mux16~5_combout ;
wire \DP|ALU|Mux16~6_combout ;
wire \DP|ALU|Mux29~6_combout ;
wire \DP|ALU|Mux28~7_combout ;
wire \DP|ALU|Mux8~8_combout ;
wire \DP|ALU|Mux10~5_combout ;
wire \DP|ALU|Mux10~6_combout ;
wire \DP|ALU|Mux9~6_combout ;
wire \DP|ALU|Mux9~7_combout ;
wire \DP|ALU|Mux30~5_combout ;
wire \DP|ALU|Mux15~6_combout ;
wire \DP|ALU|Mux15~7_combout ;
wire \DP|ALU|Mux14~6_combout ;
wire \DP|ALU|Mux14~7_combout ;
wire \DP|ALU|Mux13~5_combout ;
wire \DP|ALU|Mux13~6_combout ;
wire \DP|ALU|Mux12~5_combout ;
wire \DP|ALU|Mux12~6_combout ;
wire \DP|ALU|Mux11~5_combout ;
wire \DP|ALU|Mux11~6_combout ;
wire \DP|ALU|Mux31~12_combout ;
wire [0:0] \CC|ccif.iwait ;


memory_control CC(
	.LessThan1(LessThan1),
	.ruifdWEN_r(ruifdWEN_r),
	.ruifdREN_r(ruifdREN_r),
	.always0(always0),
	.always01(always01),
	.always02(always02),
	.ccifiwait_0(\CC|ccif.iwait[0]~0_combout ),
	.ccifiwait_01(\CC|ccif.iwait [0]),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

caches CM(
	.dpifhalt(dpifhalt),
	.ramiframload_0(ramiframload_0),
	.LessThan1(LessThan1),
	.daddr_1(daddr_1),
	.daddr_0(daddr_0),
	.daddr_3(daddr_3),
	.daddr_2(daddr_2),
	.daddr_5(daddr_5),
	.daddr_4(daddr_4),
	.daddr_7(daddr_7),
	.daddr_6(daddr_6),
	.daddr_9(daddr_9),
	.daddr_8(daddr_8),
	.daddr_11(daddr_11),
	.daddr_10(daddr_10),
	.daddr_13(daddr_13),
	.daddr_12(daddr_12),
	.daddr_15(daddr_15),
	.daddr_14(daddr_14),
	.daddr_17(daddr_17),
	.daddr_16(daddr_16),
	.daddr_19(daddr_19),
	.daddr_18(daddr_18),
	.daddr_21(daddr_21),
	.daddr_20(daddr_20),
	.daddr_23(daddr_23),
	.daddr_22(daddr_22),
	.daddr_25(daddr_25),
	.daddr_24(daddr_24),
	.daddr_27(daddr_27),
	.daddr_26(daddr_26),
	.daddr_29(daddr_29),
	.daddr_28(daddr_28),
	.daddr_31(daddr_31),
	.daddr_30(daddr_30),
	.always0(always03),
	.always1(always1),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_211),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.ccifiwait_0(\CC|ccif.iwait [0]),
	.dcifimemload_26(\CM|dcif.imemload[26]~0_combout ),
	.dcifimemload_27(\CM|dcif.imemload[27]~1_combout ),
	.dcifimemload_28(\CM|dcif.imemload[28]~2_combout ),
	.dcifimemload_29(\CM|dcif.imemload[29]~3_combout ),
	.dcifimemload_30(\CM|dcif.imemload[30]~4_combout ),
	.dcifimemload_31(\CM|dcif.imemload[31]~5_combout ),
	.dcifihit(\CM|dcif.ihit~0_combout ),
	.dcifimemload_19(\CM|dcif.imemload[19]~6_combout ),
	.dcifimemload_18(\CM|dcif.imemload[18]~7_combout ),
	.dcifimemload_16(\CM|dcif.imemload[16]~8_combout ),
	.dcifimemload_17(\CM|dcif.imemload[17]~9_combout ),
	.dcifimemload_20(dcifimemload_20),
	.dcifimemload_24(\CM|dcif.imemload[24]~11_combout ),
	.dcifimemload_23(\CM|dcif.imemload[23]~12_combout ),
	.dcifimemload_21(\CM|dcif.imemload[21]~13_combout ),
	.dcifimemload_22(\CM|dcif.imemload[22]~14_combout ),
	.dcifimemload_25(\CM|dcif.imemload[25]~15_combout ),
	.dcifimemload_3(\CM|dcif.imemload[3]~16_combout ),
	.dcifimemload_4(\CM|dcif.imemload[4]~17_combout ),
	.dcifimemload_2(\CM|dcif.imemload[2]~18_combout ),
	.dcifimemload_5(\CM|dcif.imemload[5]~19_combout ),
	.dcifimemload_0(\CM|dcif.imemload[0]~20_combout ),
	.dcifimemload_1(\CM|dcif.imemload[1]~21_combout ),
	.dcifimemload_15(\CM|dcif.imemload[15]~22_combout ),
	.dcifimemload_14(\CM|dcif.imemload[14]~23_combout ),
	.dcifimemload_13(\CM|dcif.imemload[13]~24_combout ),
	.dcifimemload_12(\CM|dcif.imemload[12]~25_combout ),
	.dcifimemload_11(\CM|dcif.imemload[11]~26_combout ),
	.dcifimemload_10(\CM|dcif.imemload[10]~27_combout ),
	.dcifimemload_9(\CM|dcif.imemload[9]~28_combout ),
	.dcifimemload_8(\CM|dcif.imemload[8]~29_combout ),
	.dcifimemload_7(\CM|dcif.imemload[7]~30_combout ),
	.dcifimemload_6(\CM|dcif.imemload[6]~31_combout ),
	.Selector0(\DP|cu|Selector0~2_combout ),
	.Mux1(\DP|ALU|Mux1~7_combout ),
	.Mux31(\DP|ALU|Mux31~0_combout ),
	.Mux11(\DP|ALU|Mux1~8_combout ),
	.Mux0(\DP|ALU|Mux0~13_combout ),
	.Mux01(\DP|ALU|Mux0~14_combout ),
	.Mux24(\DP|ALU|Mux24~9_combout ),
	.Mux25(\DP|ALU|Mux25~5_combout ),
	.Mux26(\DP|ALU|Mux26~5_combout ),
	.Mux27(\DP|ALU|Mux27~5_combout ),
	.Mux4(\DP|ALU|Mux4~6_combout ),
	.Mux5(\DP|ALU|Mux5~6_combout ),
	.Mux6(\DP|ALU|Mux6~16_combout ),
	.Mux7(\DP|ALU|Mux7~6_combout ),
	.Mux3(\DP|ALU|Mux3~7_combout ),
	.Mux2(\DP|ALU|Mux2~11_combout ),
	.Mux23(\DP|ALU|Mux23~7_combout ),
	.Mux231(\DP|ALU|Mux23~8_combout ),
	.Mux22(\DP|ALU|Mux22~5_combout ),
	.Mux221(\DP|ALU|Mux22~6_combout ),
	.Mux21(\DP|ALU|Mux21~5_combout ),
	.Mux211(\DP|ALU|Mux21~6_combout ),
	.Mux20(\DP|ALU|Mux20~5_combout ),
	.Mux201(\DP|ALU|Mux20~6_combout ),
	.Mux19(\DP|ALU|Mux19~5_combout ),
	.Mux191(\DP|ALU|Mux19~6_combout ),
	.Mux18(\DP|ALU|Mux18~8_combout ),
	.Mux181(\DP|ALU|Mux18~9_combout ),
	.Mux17(\DP|ALU|Mux17~5_combout ),
	.Mux171(\DP|ALU|Mux17~6_combout ),
	.Mux16(\DP|ALU|Mux16~5_combout ),
	.Mux161(\DP|ALU|Mux16~6_combout ),
	.Mux29(\DP|ALU|Mux29~6_combout ),
	.Mux28(\DP|ALU|Mux28~7_combout ),
	.Mux8(\DP|ALU|Mux8~8_combout ),
	.Mux10(\DP|ALU|Mux10~5_combout ),
	.Mux101(\DP|ALU|Mux10~6_combout ),
	.Mux9(\DP|ALU|Mux9~6_combout ),
	.Mux91(\DP|ALU|Mux9~7_combout ),
	.Mux30(\DP|ALU|Mux30~5_combout ),
	.Mux15(\DP|ALU|Mux15~6_combout ),
	.Mux151(\DP|ALU|Mux15~7_combout ),
	.Mux14(\DP|ALU|Mux14~6_combout ),
	.Mux141(\DP|ALU|Mux14~7_combout ),
	.Mux13(\DP|ALU|Mux13~5_combout ),
	.Mux131(\DP|ALU|Mux13~6_combout ),
	.Mux12(\DP|ALU|Mux12~5_combout ),
	.Mux121(\DP|ALU|Mux12~6_combout ),
	.Mux111(\DP|ALU|Mux11~5_combout ),
	.Mux112(\DP|ALU|Mux11~6_combout ),
	.Mux311(\DP|ALU|Mux31~12_combout ),
	.nRST(nRST),
	.CLK(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

datapath DP(
	.PC_29(PC_29),
	.PC_28(PC_28),
	.PC_31(PC_31),
	.PC_30(PC_30),
	.dpifhalt(dpifhalt),
	.PC_1(PC_1),
	.ruifdWEN_r(ruifdWEN_r),
	.ruifdREN_r(ruifdREN_r),
	.PC_0(PC_0),
	.PC_3(PC_3),
	.PC_2(PC_2),
	.PC_5(PC_5),
	.PC_4(PC_4),
	.PC_7(PC_7),
	.PC_6(PC_6),
	.PC_9(PC_9),
	.PC_8(PC_8),
	.PC_11(PC_11),
	.PC_10(PC_10),
	.PC_13(PC_13),
	.PC_12(PC_12),
	.PC_15(PC_15),
	.PC_14(PC_14),
	.PC_17(PC_17),
	.PC_16(PC_16),
	.PC_19(PC_19),
	.PC_18(PC_18),
	.PC_21(PC_21),
	.PC_20(PC_20),
	.PC_23(PC_23),
	.PC_22(PC_22),
	.PC_25(PC_25),
	.PC_24(PC_24),
	.PC_27(PC_27),
	.PC_26(PC_26),
	.ramiframload_0(ramiframload_01),
	.always1(always1),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_21),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_41),
	.ramiframload_5(ramiframload_51),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_161),
	.ramiframload_17(ramiframload_171),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_211),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_261),
	.ramiframload_27(ramiframload_271),
	.ramiframload_28(ramiframload_281),
	.ramiframload_29(ramiframload_291),
	.ramiframload_30(ramiframload_301),
	.ramiframload_31(ramiframload_311),
	.ccifiwait_0(\CC|ccif.iwait[0]~0_combout ),
	.ccifiwait_01(\CC|ccif.iwait [0]),
	.dcifimemload_26(\CM|dcif.imemload[26]~0_combout ),
	.dcifimemload_27(\CM|dcif.imemload[27]~1_combout ),
	.dcifimemload_28(\CM|dcif.imemload[28]~2_combout ),
	.dcifimemload_29(\CM|dcif.imemload[29]~3_combout ),
	.dcifimemload_30(\CM|dcif.imemload[30]~4_combout ),
	.dcifimemload_31(\CM|dcif.imemload[31]~5_combout ),
	.\dpif.ihit (\CM|dcif.ihit~0_combout ),
	.dcifimemload_19(\CM|dcif.imemload[19]~6_combout ),
	.dcifimemload_18(\CM|dcif.imemload[18]~7_combout ),
	.dcifimemload_16(\CM|dcif.imemload[16]~8_combout ),
	.dcifimemload_17(\CM|dcif.imemload[17]~9_combout ),
	.Mux63(Mux63),
	.Mux631(Mux631),
	.dcifimemload_20(dcifimemload_20),
	.dcifimemload_24(\CM|dcif.imemload[24]~11_combout ),
	.dcifimemload_23(\CM|dcif.imemload[23]~12_combout ),
	.dcifimemload_21(\CM|dcif.imemload[21]~13_combout ),
	.dcifimemload_22(\CM|dcif.imemload[22]~14_combout ),
	.dcifimemload_25(\CM|dcif.imemload[25]~15_combout ),
	.dcifimemload_3(\CM|dcif.imemload[3]~16_combout ),
	.dcifimemload_4(\CM|dcif.imemload[4]~17_combout ),
	.dcifimemload_2(\CM|dcif.imemload[2]~18_combout ),
	.dcifimemload_5(\CM|dcif.imemload[5]~19_combout ),
	.dcifimemload_0(\CM|dcif.imemload[0]~20_combout ),
	.dcifimemload_1(\CM|dcif.imemload[1]~21_combout ),
	.Mux33(Mux33),
	.dcifimemload_15(\CM|dcif.imemload[15]~22_combout ),
	.Mux331(Mux331),
	.Mux34(Mux34),
	.Mux341(Mux341),
	.Mux35(Mux35),
	.Mux351(Mux351),
	.Mux36(Mux36),
	.Mux361(Mux361),
	.Mux37(Mux37),
	.Mux371(Mux371),
	.Mux38(Mux38),
	.Mux381(Mux381),
	.Mux39(Mux39),
	.Mux391(Mux391),
	.Mux40(Mux40),
	.Mux401(Mux401),
	.Mux41(Mux41),
	.Mux411(Mux411),
	.Mux42(Mux42),
	.Mux421(Mux421),
	.Mux43(Mux43),
	.Mux431(Mux431),
	.Mux44(Mux44),
	.Mux441(Mux441),
	.Mux45(Mux45),
	.Mux451(Mux451),
	.Mux46(Mux46),
	.Mux461(Mux461),
	.Mux47(Mux47),
	.Mux471(Mux471),
	.Mux48(Mux48),
	.Mux481(Mux481),
	.Mux49(Mux49),
	.Mux491(Mux491),
	.dcifimemload_14(\CM|dcif.imemload[14]~23_combout ),
	.Mux50(Mux50),
	.Mux501(Mux501),
	.dcifimemload_13(\CM|dcif.imemload[13]~24_combout ),
	.Mux51(Mux51),
	.Mux511(Mux511),
	.dcifimemload_12(\CM|dcif.imemload[12]~25_combout ),
	.Mux52(Mux52),
	.Mux521(Mux521),
	.dcifimemload_11(\CM|dcif.imemload[11]~26_combout ),
	.Mux53(Mux53),
	.Mux531(Mux531),
	.dcifimemload_10(\CM|dcif.imemload[10]~27_combout ),
	.Mux54(Mux54),
	.Mux541(Mux541),
	.dcifimemload_9(\CM|dcif.imemload[9]~28_combout ),
	.Mux55(Mux55),
	.Mux551(Mux551),
	.dcifimemload_8(\CM|dcif.imemload[8]~29_combout ),
	.Mux56(Mux56),
	.Mux561(Mux561),
	.dcifimemload_7(\CM|dcif.imemload[7]~30_combout ),
	.Mux57(Mux57),
	.Mux571(Mux571),
	.dcifimemload_6(\CM|dcif.imemload[6]~31_combout ),
	.Mux58(Mux58),
	.Mux581(Mux581),
	.Mux59(Mux59),
	.Mux591(Mux591),
	.Mux60(Mux60),
	.Mux601(Mux601),
	.Mux61(Mux61),
	.Mux611(Mux611),
	.Mux62(Mux62),
	.Mux621(Mux621),
	.Mux32(Mux32),
	.Mux321(Mux321),
	.Selector0(\DP|cu|Selector0~2_combout ),
	.Mux1(\DP|ALU|Mux1~7_combout ),
	.Mux31(\DP|ALU|Mux31~0_combout ),
	.Mux11(\DP|ALU|Mux1~8_combout ),
	.Mux0(\DP|ALU|Mux0~13_combout ),
	.Mux01(\DP|ALU|Mux0~14_combout ),
	.Mux24(\DP|ALU|Mux24~9_combout ),
	.Mux25(\DP|ALU|Mux25~5_combout ),
	.Mux26(\DP|ALU|Mux26~5_combout ),
	.Mux27(\DP|ALU|Mux27~5_combout ),
	.Mux4(\DP|ALU|Mux4~6_combout ),
	.Mux5(\DP|ALU|Mux5~6_combout ),
	.Mux6(\DP|ALU|Mux6~16_combout ),
	.Mux7(\DP|ALU|Mux7~6_combout ),
	.Mux3(\DP|ALU|Mux3~7_combout ),
	.Mux2(\DP|ALU|Mux2~11_combout ),
	.Mux23(\DP|ALU|Mux23~7_combout ),
	.Mux231(\DP|ALU|Mux23~8_combout ),
	.Mux22(\DP|ALU|Mux22~5_combout ),
	.Mux221(\DP|ALU|Mux22~6_combout ),
	.Mux21(\DP|ALU|Mux21~5_combout ),
	.Mux211(\DP|ALU|Mux21~6_combout ),
	.Mux20(\DP|ALU|Mux20~5_combout ),
	.Mux201(\DP|ALU|Mux20~6_combout ),
	.Mux19(\DP|ALU|Mux19~5_combout ),
	.Mux191(\DP|ALU|Mux19~6_combout ),
	.Mux18(\DP|ALU|Mux18~8_combout ),
	.Mux181(\DP|ALU|Mux18~9_combout ),
	.Mux17(\DP|ALU|Mux17~5_combout ),
	.Mux171(\DP|ALU|Mux17~6_combout ),
	.Mux16(\DP|ALU|Mux16~5_combout ),
	.Mux161(\DP|ALU|Mux16~6_combout ),
	.Mux29(\DP|ALU|Mux29~6_combout ),
	.Mux28(\DP|ALU|Mux28~7_combout ),
	.Mux8(\DP|ALU|Mux8~8_combout ),
	.Mux10(\DP|ALU|Mux10~5_combout ),
	.Mux101(\DP|ALU|Mux10~6_combout ),
	.Mux9(\DP|ALU|Mux9~6_combout ),
	.Mux91(\DP|ALU|Mux9~7_combout ),
	.Mux30(\DP|ALU|Mux30~5_combout ),
	.Mux15(\DP|ALU|Mux15~6_combout ),
	.Mux151(\DP|ALU|Mux15~7_combout ),
	.Mux14(\DP|ALU|Mux14~6_combout ),
	.Mux141(\DP|ALU|Mux14~7_combout ),
	.Mux13(\DP|ALU|Mux13~5_combout ),
	.Mux131(\DP|ALU|Mux13~6_combout ),
	.Mux12(\DP|ALU|Mux12~5_combout ),
	.Mux121(\DP|ALU|Mux12~6_combout ),
	.Mux111(\DP|ALU|Mux11~5_combout ),
	.Mux112(\DP|ALU|Mux11~6_combout ),
	.Mux311(\DP|ALU|Mux31~12_combout ),
	.CLK(CLK),
	.nRST(nRST1),
	.dpifhalt1(dpifhalt1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module caches (
	dpifhalt,
	ramiframload_0,
	LessThan1,
	daddr_1,
	daddr_0,
	daddr_3,
	daddr_2,
	daddr_5,
	daddr_4,
	daddr_7,
	daddr_6,
	daddr_9,
	daddr_8,
	daddr_11,
	daddr_10,
	daddr_13,
	daddr_12,
	daddr_15,
	daddr_14,
	daddr_17,
	daddr_16,
	daddr_19,
	daddr_18,
	daddr_21,
	daddr_20,
	daddr_23,
	daddr_22,
	daddr_25,
	daddr_24,
	daddr_27,
	daddr_26,
	daddr_29,
	daddr_28,
	daddr_31,
	daddr_30,
	always0,
	always1,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ccifiwait_0,
	dcifimemload_26,
	dcifimemload_27,
	dcifimemload_28,
	dcifimemload_29,
	dcifimemload_30,
	dcifimemload_31,
	dcifihit,
	dcifimemload_19,
	dcifimemload_18,
	dcifimemload_16,
	dcifimemload_17,
	dcifimemload_20,
	dcifimemload_24,
	dcifimemload_23,
	dcifimemload_21,
	dcifimemload_22,
	dcifimemload_25,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_0,
	dcifimemload_1,
	dcifimemload_15,
	dcifimemload_14,
	dcifimemload_13,
	dcifimemload_12,
	dcifimemload_11,
	dcifimemload_10,
	dcifimemload_9,
	dcifimemload_8,
	dcifimemload_7,
	dcifimemload_6,
	Selector0,
	Mux1,
	Mux31,
	Mux11,
	Mux0,
	Mux01,
	Mux24,
	Mux25,
	Mux26,
	Mux27,
	Mux4,
	Mux5,
	Mux6,
	Mux7,
	Mux3,
	Mux2,
	Mux23,
	Mux231,
	Mux22,
	Mux221,
	Mux21,
	Mux211,
	Mux20,
	Mux201,
	Mux19,
	Mux191,
	Mux18,
	Mux181,
	Mux17,
	Mux171,
	Mux16,
	Mux161,
	Mux29,
	Mux28,
	Mux8,
	Mux10,
	Mux101,
	Mux9,
	Mux91,
	Mux30,
	Mux15,
	Mux151,
	Mux14,
	Mux141,
	Mux13,
	Mux131,
	Mux12,
	Mux121,
	Mux111,
	Mux112,
	Mux311,
	nRST,
	CLK,
	devpor,
	devclrn,
	devoe);
input 	dpifhalt;
input 	ramiframload_0;
input 	LessThan1;
output 	daddr_1;
output 	daddr_0;
output 	daddr_3;
output 	daddr_2;
output 	daddr_5;
output 	daddr_4;
output 	daddr_7;
output 	daddr_6;
output 	daddr_9;
output 	daddr_8;
output 	daddr_11;
output 	daddr_10;
output 	daddr_13;
output 	daddr_12;
output 	daddr_15;
output 	daddr_14;
output 	daddr_17;
output 	daddr_16;
output 	daddr_19;
output 	daddr_18;
output 	daddr_21;
output 	daddr_20;
output 	daddr_23;
output 	daddr_22;
output 	daddr_25;
output 	daddr_24;
output 	daddr_27;
output 	daddr_26;
output 	daddr_29;
output 	daddr_28;
output 	daddr_31;
output 	daddr_30;
input 	always0;
input 	always1;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	ccifiwait_0;
output 	dcifimemload_26;
output 	dcifimemload_27;
output 	dcifimemload_28;
output 	dcifimemload_29;
output 	dcifimemload_30;
output 	dcifimemload_31;
output 	dcifihit;
output 	dcifimemload_19;
output 	dcifimemload_18;
output 	dcifimemload_16;
output 	dcifimemload_17;
output 	dcifimemload_20;
output 	dcifimemload_24;
output 	dcifimemload_23;
output 	dcifimemload_21;
output 	dcifimemload_22;
output 	dcifimemload_25;
output 	dcifimemload_3;
output 	dcifimemload_4;
output 	dcifimemload_2;
output 	dcifimemload_5;
output 	dcifimemload_0;
output 	dcifimemload_1;
output 	dcifimemload_15;
output 	dcifimemload_14;
output 	dcifimemload_13;
output 	dcifimemload_12;
output 	dcifimemload_11;
output 	dcifimemload_10;
output 	dcifimemload_9;
output 	dcifimemload_8;
output 	dcifimemload_7;
output 	dcifimemload_6;
input 	Selector0;
input 	Mux1;
input 	Mux31;
input 	Mux11;
input 	Mux0;
input 	Mux01;
input 	Mux24;
input 	Mux25;
input 	Mux26;
input 	Mux27;
input 	Mux4;
input 	Mux5;
input 	Mux6;
input 	Mux7;
input 	Mux3;
input 	Mux2;
input 	Mux23;
input 	Mux231;
input 	Mux22;
input 	Mux221;
input 	Mux21;
input 	Mux211;
input 	Mux20;
input 	Mux201;
input 	Mux19;
input 	Mux191;
input 	Mux18;
input 	Mux181;
input 	Mux17;
input 	Mux171;
input 	Mux16;
input 	Mux161;
input 	Mux29;
input 	Mux28;
input 	Mux8;
input 	Mux10;
input 	Mux101;
input 	Mux9;
input 	Mux91;
input 	Mux30;
input 	Mux15;
input 	Mux151;
input 	Mux14;
input 	Mux141;
input 	Mux13;
input 	Mux131;
input 	Mux12;
input 	Mux121;
input 	Mux111;
input 	Mux112;
input 	Mux311;
input 	nRST;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \daddr~0_combout ;
wire \instr[1]~0_combout ;
wire \daddr~1_combout ;
wire \daddr~2_combout ;
wire \daddr~3_combout ;
wire \daddr~4_combout ;
wire \daddr~5_combout ;
wire \daddr~6_combout ;
wire \daddr~7_combout ;
wire \daddr~8_combout ;
wire \daddr~9_combout ;
wire \daddr~10_combout ;
wire \daddr~11_combout ;
wire \daddr~12_combout ;
wire \daddr~13_combout ;
wire \daddr~14_combout ;
wire \daddr~15_combout ;
wire \daddr~16_combout ;
wire \daddr~17_combout ;
wire \daddr~18_combout ;
wire \daddr~19_combout ;
wire \daddr~20_combout ;
wire \daddr~21_combout ;
wire \daddr~22_combout ;
wire \daddr~23_combout ;
wire \daddr~24_combout ;
wire \daddr~25_combout ;
wire \daddr~26_combout ;
wire \daddr~27_combout ;
wire \daddr~28_combout ;
wire \daddr~29_combout ;
wire \daddr~30_combout ;
wire \daddr~31_combout ;
wire \instr~1_combout ;
wire \instr~2_combout ;
wire \instr~3_combout ;
wire \instr~4_combout ;
wire \instr~5_combout ;
wire \instr~6_combout ;
wire \instr~7_combout ;
wire \instr~8_combout ;
wire \instr~9_combout ;
wire \instr~10_combout ;
wire \instr~11_combout ;
wire \instr~12_combout ;
wire \instr~13_combout ;
wire \instr~14_combout ;
wire \instr~15_combout ;
wire \instr~16_combout ;
wire \instr~17_combout ;
wire \instr~18_combout ;
wire \instr~19_combout ;
wire \instr~20_combout ;
wire \instr~21_combout ;
wire \instr~22_combout ;
wire \instr~23_combout ;
wire \instr~24_combout ;
wire \instr~25_combout ;
wire \instr~26_combout ;
wire \instr~27_combout ;
wire \instr~28_combout ;
wire \instr~29_combout ;
wire \instr~30_combout ;
wire \instr~31_combout ;
wire \instr~32_combout ;
wire [31:0] instr;


// Location: FF_X55_Y34_N17
dffeas \daddr[1] (
	.clk(CLK),
	.d(\daddr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_1),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[1] .is_wysiwyg = "true";
defparam \daddr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N9
dffeas \daddr[0] (
	.clk(CLK),
	.d(\daddr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_0),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[0] .is_wysiwyg = "true";
defparam \daddr[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N13
dffeas \daddr[3] (
	.clk(CLK),
	.d(\daddr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_3),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[3] .is_wysiwyg = "true";
defparam \daddr[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N29
dffeas \daddr[2] (
	.clk(CLK),
	.d(\daddr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_2),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[2] .is_wysiwyg = "true";
defparam \daddr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N15
dffeas \daddr[5] (
	.clk(CLK),
	.d(\daddr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_5),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[5] .is_wysiwyg = "true";
defparam \daddr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N25
dffeas \daddr[4] (
	.clk(CLK),
	.d(\daddr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_4),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[4] .is_wysiwyg = "true";
defparam \daddr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y44_N5
dffeas \daddr[7] (
	.clk(CLK),
	.d(\daddr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_7),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[7] .is_wysiwyg = "true";
defparam \daddr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N19
dffeas \daddr[6] (
	.clk(CLK),
	.d(\daddr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_6),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[6] .is_wysiwyg = "true";
defparam \daddr[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N29
dffeas \daddr[9] (
	.clk(CLK),
	.d(\daddr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_9),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[9] .is_wysiwyg = "true";
defparam \daddr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N31
dffeas \daddr[8] (
	.clk(CLK),
	.d(\daddr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_8),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[8] .is_wysiwyg = "true";
defparam \daddr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N17
dffeas \daddr[11] (
	.clk(CLK),
	.d(\daddr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_11),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[11] .is_wysiwyg = "true";
defparam \daddr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N9
dffeas \daddr[10] (
	.clk(CLK),
	.d(\daddr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_10),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[10] .is_wysiwyg = "true";
defparam \daddr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y43_N21
dffeas \daddr[13] (
	.clk(CLK),
	.d(\daddr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_13),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[13] .is_wysiwyg = "true";
defparam \daddr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N21
dffeas \daddr[12] (
	.clk(CLK),
	.d(\daddr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_12),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[12] .is_wysiwyg = "true";
defparam \daddr[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N7
dffeas \daddr[15] (
	.clk(CLK),
	.d(\daddr~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_15),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[15] .is_wysiwyg = "true";
defparam \daddr[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N17
dffeas \daddr[14] (
	.clk(CLK),
	.d(\daddr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_14),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[14] .is_wysiwyg = "true";
defparam \daddr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N5
dffeas \daddr[17] (
	.clk(CLK),
	.d(\daddr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_17),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[17] .is_wysiwyg = "true";
defparam \daddr[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N23
dffeas \daddr[16] (
	.clk(CLK),
	.d(\daddr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_16),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[16] .is_wysiwyg = "true";
defparam \daddr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y43_N15
dffeas \daddr[19] (
	.clk(CLK),
	.d(\daddr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_19),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[19] .is_wysiwyg = "true";
defparam \daddr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N27
dffeas \daddr[18] (
	.clk(CLK),
	.d(\daddr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_18),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[18] .is_wysiwyg = "true";
defparam \daddr[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N17
dffeas \daddr[21] (
	.clk(CLK),
	.d(\daddr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_21),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[21] .is_wysiwyg = "true";
defparam \daddr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y43_N25
dffeas \daddr[20] (
	.clk(CLK),
	.d(\daddr~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_20),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[20] .is_wysiwyg = "true";
defparam \daddr[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N21
dffeas \daddr[23] (
	.clk(CLK),
	.d(\daddr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_23),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[23] .is_wysiwyg = "true";
defparam \daddr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N11
dffeas \daddr[22] (
	.clk(CLK),
	.d(\daddr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_22),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[22] .is_wysiwyg = "true";
defparam \daddr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N5
dffeas \daddr[25] (
	.clk(CLK),
	.d(\daddr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_25),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[25] .is_wysiwyg = "true";
defparam \daddr[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y42_N17
dffeas \daddr[24] (
	.clk(CLK),
	.d(\daddr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_24),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[24] .is_wysiwyg = "true";
defparam \daddr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N7
dffeas \daddr[27] (
	.clk(CLK),
	.d(\daddr~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_27),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[27] .is_wysiwyg = "true";
defparam \daddr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N3
dffeas \daddr[26] (
	.clk(CLK),
	.d(\daddr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_26),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[26] .is_wysiwyg = "true";
defparam \daddr[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N9
dffeas \daddr[29] (
	.clk(CLK),
	.d(\daddr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_29),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[29] .is_wysiwyg = "true";
defparam \daddr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N31
dffeas \daddr[28] (
	.clk(CLK),
	.d(\daddr~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_28),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[28] .is_wysiwyg = "true";
defparam \daddr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N5
dffeas \daddr[31] (
	.clk(CLK),
	.d(\daddr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_31),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[31] .is_wysiwyg = "true";
defparam \daddr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N25
dffeas \daddr[30] (
	.clk(CLK),
	.d(\daddr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_30),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[30] .is_wysiwyg = "true";
defparam \daddr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N2
cycloneive_lcell_comb \dcif.imemload[26]~0 (
// Equation(s):
// dcifimemload_26 = (ccifiwait_01 & (((instr[26])))) # (!ccifiwait_01 & (ramiframload_26 & ((always1))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_26),
	.datac(instr[26]),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_26),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[26]~0 .lut_mask = 16'hE4A0;
defparam \dcif.imemload[26]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N28
cycloneive_lcell_comb \dcif.imemload[27]~1 (
// Equation(s):
// dcifimemload_27 = (ccifiwait_01 & (((instr[27])))) # (!ccifiwait_01 & ((ramiframload_27) # ((!always1))))

	.dataa(ramiframload_27),
	.datab(always1),
	.datac(instr[27]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_27),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[27]~1 .lut_mask = 16'hF0BB;
defparam \dcif.imemload[27]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N14
cycloneive_lcell_comb \dcif.imemload[28]~2 (
// Equation(s):
// dcifimemload_28 = (ccifiwait_01 & (((instr[28])))) # (!ccifiwait_01 & (((ramiframload_28)) # (!always1)))

	.dataa(ccifiwait_0),
	.datab(always1),
	.datac(instr[28]),
	.datad(ramiframload_28),
	.cin(gnd),
	.combout(dcifimemload_28),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[28]~2 .lut_mask = 16'hF5B1;
defparam \dcif.imemload[28]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N8
cycloneive_lcell_comb \dcif.imemload[29]~3 (
// Equation(s):
// dcifimemload_29 = (ccifiwait_01 & (((instr[29])))) # (!ccifiwait_01 & ((ramiframload_29) # ((!always1))))

	.dataa(ramiframload_29),
	.datab(always1),
	.datac(instr[29]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_29),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[29]~3 .lut_mask = 16'hF0BB;
defparam \dcif.imemload[29]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N18
cycloneive_lcell_comb \dcif.imemload[30]~4 (
// Equation(s):
// dcifimemload_30 = (ccifiwait_01 & (((instr[30])))) # (!ccifiwait_01 & (ramiframload_30 & (always1)))

	.dataa(ramiframload_30),
	.datab(always1),
	.datac(instr[30]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_30),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[30]~4 .lut_mask = 16'hF088;
defparam \dcif.imemload[30]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N4
cycloneive_lcell_comb \dcif.imemload[31]~5 (
// Equation(s):
// dcifimemload_31 = (ccifiwait_01 & (((instr[31])))) # (!ccifiwait_01 & ((ramiframload_31) # ((!always1))))

	.dataa(ramiframload_31),
	.datab(always1),
	.datac(instr[31]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_31),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[31]~5 .lut_mask = 16'hF0BB;
defparam \dcif.imemload[31]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N4
cycloneive_lcell_comb \dcif.ihit~0 (
// Equation(s):
// dcifihit = (!dpifhalt & !ccifiwait_01)

	.dataa(gnd),
	.datab(dpifhalt),
	.datac(gnd),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifihit),
	.cout());
// synopsys translate_off
defparam \dcif.ihit~0 .lut_mask = 16'h0033;
defparam \dcif.ihit~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N30
cycloneive_lcell_comb \dcif.imemload[19]~6 (
// Equation(s):
// dcifimemload_19 = (ccifiwait_01 & (instr[19])) # (!ccifiwait_01 & ((ramiframload_19)))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(instr[19]),
	.datad(ramiframload_19),
	.cin(gnd),
	.combout(dcifimemload_19),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[19]~6 .lut_mask = 16'hF5A0;
defparam \dcif.imemload[19]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N26
cycloneive_lcell_comb \dcif.imemload[18]~7 (
// Equation(s):
// dcifimemload_18 = (ccifiwait_01 & (instr[18])) # (!ccifiwait_01 & ((ramiframload_18)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[18]),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(dcifimemload_18),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[18]~7 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[18]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N4
cycloneive_lcell_comb \dcif.imemload[16]~8 (
// Equation(s):
// dcifimemload_16 = (ccifiwait_01 & (((instr[16])))) # (!ccifiwait_01 & (((ramiframload_16)) # (!always1)))

	.dataa(always1),
	.datab(ccifiwait_0),
	.datac(instr[16]),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(dcifimemload_16),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[16]~8 .lut_mask = 16'hF3D1;
defparam \dcif.imemload[16]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N14
cycloneive_lcell_comb \dcif.imemload[17]~9 (
// Equation(s):
// dcifimemload_17 = (ccifiwait_01 & (((instr[17])))) # (!ccifiwait_01 & (always1 & ((ramiframload_17))))

	.dataa(always1),
	.datab(ccifiwait_0),
	.datac(instr[17]),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(dcifimemload_17),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[17]~9 .lut_mask = 16'hE2C0;
defparam \dcif.imemload[17]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N12
cycloneive_lcell_comb \dcif.imemload[20]~10 (
// Equation(s):
// dcifimemload_20 = (ccifiwait_01 & (instr[20])) # (!ccifiwait_01 & ((ramiframload_20)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[20]),
	.datad(ramiframload_20),
	.cin(gnd),
	.combout(dcifimemload_20),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[20]~10 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[20]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N26
cycloneive_lcell_comb \dcif.imemload[24]~11 (
// Equation(s):
// dcifimemload_24 = (ccifiwait_01 & (instr[24])) # (!ccifiwait_01 & ((ramiframload_24)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[24]),
	.datad(ramiframload_24),
	.cin(gnd),
	.combout(dcifimemload_24),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[24]~11 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[24]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N12
cycloneive_lcell_comb \dcif.imemload[23]~12 (
// Equation(s):
// dcifimemload_23 = (ccifiwait_01 & (instr[23])) # (!ccifiwait_01 & ((ramiframload_23)))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(instr[23]),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(dcifimemload_23),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[23]~12 .lut_mask = 16'hF5A0;
defparam \dcif.imemload[23]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N4
cycloneive_lcell_comb \dcif.imemload[21]~13 (
// Equation(s):
// dcifimemload_21 = (ccifiwait_01 & (instr[21])) # (!ccifiwait_01 & ((ramiframload_211)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[21]),
	.datad(ramiframload_21),
	.cin(gnd),
	.combout(dcifimemload_21),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[21]~13 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[21]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N16
cycloneive_lcell_comb \dcif.imemload[22]~14 (
// Equation(s):
// dcifimemload_22 = (ccifiwait_01 & (instr[22])) # (!ccifiwait_01 & ((ramiframload_22)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[22]),
	.datad(ramiframload_22),
	.cin(gnd),
	.combout(dcifimemload_22),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[22]~14 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[22]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N20
cycloneive_lcell_comb \dcif.imemload[25]~15 (
// Equation(s):
// dcifimemload_25 = (ccifiwait_01 & (instr[25])) # (!ccifiwait_01 & ((ramiframload_25)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[25]),
	.datad(ramiframload_25),
	.cin(gnd),
	.combout(dcifimemload_25),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[25]~15 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[25]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N30
cycloneive_lcell_comb \dcif.imemload[3]~16 (
// Equation(s):
// dcifimemload_3 = (ccifiwait_01 & (instr[3])) # (!ccifiwait_01 & ((ramiframload_3)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[3]),
	.datad(ramiframload_3),
	.cin(gnd),
	.combout(dcifimemload_3),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[3]~16 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[3]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N4
cycloneive_lcell_comb \dcif.imemload[4]~17 (
// Equation(s):
// dcifimemload_4 = (ccifiwait_01 & (((instr[4])))) # (!ccifiwait_01 & (((ramiframload_4)) # (!always1)))

	.dataa(always1),
	.datab(ccifiwait_0),
	.datac(instr[4]),
	.datad(ramiframload_4),
	.cin(gnd),
	.combout(dcifimemload_4),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[4]~17 .lut_mask = 16'hF3D1;
defparam \dcif.imemload[4]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N22
cycloneive_lcell_comb \dcif.imemload[2]~18 (
// Equation(s):
// dcifimemload_2 = (ccifiwait_01 & (((instr[2])))) # (!ccifiwait_01 & (always1 & ((ramiframload_2))))

	.dataa(always1),
	.datab(ccifiwait_0),
	.datac(instr[2]),
	.datad(ramiframload_2),
	.cin(gnd),
	.combout(dcifimemload_2),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[2]~18 .lut_mask = 16'hE2C0;
defparam \dcif.imemload[2]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N20
cycloneive_lcell_comb \dcif.imemload[5]~19 (
// Equation(s):
// dcifimemload_5 = (ccifiwait_01 & (((instr[5])))) # (!ccifiwait_01 & (always1 & ((ramiframload_5))))

	.dataa(always1),
	.datab(ccifiwait_0),
	.datac(instr[5]),
	.datad(ramiframload_5),
	.cin(gnd),
	.combout(dcifimemload_5),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[5]~19 .lut_mask = 16'hE2C0;
defparam \dcif.imemload[5]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N10
cycloneive_lcell_comb \dcif.imemload[0]~20 (
// Equation(s):
// dcifimemload_0 = (ccifiwait_01 & (((instr[0])))) # (!ccifiwait_01 & (((ramiframload_0)) # (!always1)))

	.dataa(always1),
	.datab(ccifiwait_0),
	.datac(instr[0]),
	.datad(ramiframload_0),
	.cin(gnd),
	.combout(dcifimemload_0),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[0]~20 .lut_mask = 16'hF3D1;
defparam \dcif.imemload[0]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N14
cycloneive_lcell_comb \dcif.imemload[1]~21 (
// Equation(s):
// dcifimemload_1 = (ccifiwait_01 & (instr[1])) # (!ccifiwait_01 & ((ramiframload_1)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[1]),
	.datad(ramiframload_1),
	.cin(gnd),
	.combout(dcifimemload_1),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[1]~21 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[1]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N24
cycloneive_lcell_comb \dcif.imemload[15]~22 (
// Equation(s):
// dcifimemload_15 = (ccifiwait_01 & ((instr[15]))) # (!ccifiwait_01 & (ramiframload_15))

	.dataa(ramiframload_15),
	.datab(gnd),
	.datac(instr[15]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_15),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[15]~22 .lut_mask = 16'hF0AA;
defparam \dcif.imemload[15]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N28
cycloneive_lcell_comb \dcif.imemload[14]~23 (
// Equation(s):
// dcifimemload_14 = (ccifiwait_01 & ((instr[14]))) # (!ccifiwait_01 & (ramiframload_14))

	.dataa(ramiframload_14),
	.datab(gnd),
	.datac(instr[14]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_14),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[14]~23 .lut_mask = 16'hF0AA;
defparam \dcif.imemload[14]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N6
cycloneive_lcell_comb \dcif.imemload[13]~24 (
// Equation(s):
// dcifimemload_13 = (ccifiwait_01 & (instr[13])) # (!ccifiwait_01 & ((ramiframload_13)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[13]),
	.datad(ramiframload_13),
	.cin(gnd),
	.combout(dcifimemload_13),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[13]~24 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[13]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N4
cycloneive_lcell_comb \dcif.imemload[12]~25 (
// Equation(s):
// dcifimemload_12 = (ccifiwait_01 & (instr[12])) # (!ccifiwait_01 & ((ramiframload_12)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[12]),
	.datad(ramiframload_12),
	.cin(gnd),
	.combout(dcifimemload_12),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[12]~25 .lut_mask = 16'hF3C0;
defparam \dcif.imemload[12]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N18
cycloneive_lcell_comb \dcif.imemload[11]~26 (
// Equation(s):
// dcifimemload_11 = (ccifiwait_01 & ((instr[11]))) # (!ccifiwait_01 & (ramiframload_11))

	.dataa(gnd),
	.datab(ramiframload_11),
	.datac(instr[11]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_11),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[11]~26 .lut_mask = 16'hF0CC;
defparam \dcif.imemload[11]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N8
cycloneive_lcell_comb \dcif.imemload[10]~27 (
// Equation(s):
// dcifimemload_10 = (ccifiwait_01 & ((instr[10]))) # (!ccifiwait_01 & (ramiframload_10))

	.dataa(gnd),
	.datab(ramiframload_10),
	.datac(instr[10]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_10),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[10]~27 .lut_mask = 16'hF0CC;
defparam \dcif.imemload[10]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N26
cycloneive_lcell_comb \dcif.imemload[9]~28 (
// Equation(s):
// dcifimemload_9 = (ccifiwait_01 & ((instr[9]))) # (!ccifiwait_01 & (ramiframload_9))

	.dataa(gnd),
	.datab(ramiframload_9),
	.datac(instr[9]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_9),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[9]~28 .lut_mask = 16'hF0CC;
defparam \dcif.imemload[9]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N4
cycloneive_lcell_comb \dcif.imemload[8]~29 (
// Equation(s):
// dcifimemload_8 = (ccifiwait_01 & ((instr[8]))) # (!ccifiwait_01 & (ramiframload_8))

	.dataa(ramiframload_8),
	.datab(gnd),
	.datac(instr[8]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_8),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[8]~29 .lut_mask = 16'hF0AA;
defparam \dcif.imemload[8]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N22
cycloneive_lcell_comb \dcif.imemload[7]~30 (
// Equation(s):
// dcifimemload_7 = (ccifiwait_01 & ((instr[7]))) # (!ccifiwait_01 & (ramiframload_7))

	.dataa(gnd),
	.datab(ramiframload_7),
	.datac(instr[7]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_7),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[7]~30 .lut_mask = 16'hF0CC;
defparam \dcif.imemload[7]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N20
cycloneive_lcell_comb \dcif.imemload[6]~31 (
// Equation(s):
// dcifimemload_6 = (ccifiwait_01 & (instr[6])) # (!ccifiwait_01 & ((ramiframload_6)))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(instr[6]),
	.datad(ramiframload_6),
	.cin(gnd),
	.combout(dcifimemload_6),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[6]~31 .lut_mask = 16'hF5A0;
defparam \dcif.imemload[6]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N16
cycloneive_lcell_comb \daddr~0 (
// Equation(s):
// \daddr~0_combout  = (\nRST~input_o  & Mux301)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Mux30),
	.cin(gnd),
	.combout(\daddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~0 .lut_mask = 16'hF000;
defparam \daddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N12
cycloneive_lcell_comb \instr[1]~0 (
// Equation(s):
// \instr[1]~0_combout  = ((!ccifiwait_01 & !dpifhalt)) # (!\nRST~input_o )

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(nRST),
	.datad(dpifhalt),
	.cin(gnd),
	.combout(\instr[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \instr[1]~0 .lut_mask = 16'h0F5F;
defparam \instr[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N8
cycloneive_lcell_comb \daddr~1 (
// Equation(s):
// \daddr~1_combout  = (Mux312 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux311),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~1 .lut_mask = 16'hF000;
defparam \daddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N12
cycloneive_lcell_comb \daddr~2 (
// Equation(s):
// \daddr~2_combout  = (Mux281 & \nRST~input_o )

	.dataa(gnd),
	.datab(Mux28),
	.datac(nRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~2 .lut_mask = 16'hC0C0;
defparam \daddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N28
cycloneive_lcell_comb \daddr~3 (
// Equation(s):
// \daddr~3_combout  = (\nRST~input_o  & Mux291)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Mux29),
	.cin(gnd),
	.combout(\daddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~3 .lut_mask = 16'hF000;
defparam \daddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N14
cycloneive_lcell_comb \daddr~4 (
// Equation(s):
// \daddr~4_combout  = (!Selector0 & (\nRST~input_o  & Mux261))

	.dataa(Selector0),
	.datab(nRST),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\daddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~4 .lut_mask = 16'h4400;
defparam \daddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N24
cycloneive_lcell_comb \daddr~5 (
// Equation(s):
// \daddr~5_combout  = (!Selector0 & (\nRST~input_o  & Mux271))

	.dataa(Selector0),
	.datab(gnd),
	.datac(nRST),
	.datad(Mux27),
	.cin(gnd),
	.combout(\daddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~5 .lut_mask = 16'h5000;
defparam \daddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N4
cycloneive_lcell_comb \daddr~6 (
// Equation(s):
// \daddr~6_combout  = (\nRST~input_o  & (Mux241 & !Selector0))

	.dataa(nRST),
	.datab(gnd),
	.datac(Mux24),
	.datad(Selector0),
	.cin(gnd),
	.combout(\daddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~6 .lut_mask = 16'h00A0;
defparam \daddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N18
cycloneive_lcell_comb \daddr~7 (
// Equation(s):
// \daddr~7_combout  = (Mux251 & (\nRST~input_o  & !Selector0))

	.dataa(gnd),
	.datab(Mux25),
	.datac(nRST),
	.datad(Selector0),
	.cin(gnd),
	.combout(\daddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~7 .lut_mask = 16'h00C0;
defparam \daddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N28
cycloneive_lcell_comb \daddr~8 (
// Equation(s):
// \daddr~8_combout  = (\nRST~input_o  & ((Mux221) # ((Mux222 & Mux311))))

	.dataa(nRST),
	.datab(Mux221),
	.datac(Mux31),
	.datad(Mux22),
	.cin(gnd),
	.combout(\daddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~8 .lut_mask = 16'hAA80;
defparam \daddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N30
cycloneive_lcell_comb \daddr~9 (
// Equation(s):
// \daddr~9_combout  = (\nRST~input_o  & ((Mux231) # ((Mux232 & Mux311))))

	.dataa(nRST),
	.datab(Mux231),
	.datac(Mux31),
	.datad(Mux23),
	.cin(gnd),
	.combout(\daddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~9 .lut_mask = 16'hAA80;
defparam \daddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N16
cycloneive_lcell_comb \daddr~10 (
// Equation(s):
// \daddr~10_combout  = (\nRST~input_o  & ((Mux201) # ((Mux311 & Mux202))))

	.dataa(Mux31),
	.datab(nRST),
	.datac(Mux201),
	.datad(Mux20),
	.cin(gnd),
	.combout(\daddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~10 .lut_mask = 16'hCC80;
defparam \daddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N8
cycloneive_lcell_comb \daddr~11 (
// Equation(s):
// \daddr~11_combout  = (\nRST~input_o  & ((Mux211) # ((Mux311 & Mux212))))

	.dataa(nRST),
	.datab(Mux31),
	.datac(Mux21),
	.datad(Mux211),
	.cin(gnd),
	.combout(\daddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~11 .lut_mask = 16'hA8A0;
defparam \daddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N20
cycloneive_lcell_comb \daddr~12 (
// Equation(s):
// \daddr~12_combout  = (\nRST~input_o  & ((Mux181) # ((Mux311 & Mux182))))

	.dataa(Mux18),
	.datab(Mux31),
	.datac(nRST),
	.datad(Mux181),
	.cin(gnd),
	.combout(\daddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~12 .lut_mask = 16'hE0A0;
defparam \daddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N20
cycloneive_lcell_comb \daddr~13 (
// Equation(s):
// \daddr~13_combout  = (\nRST~input_o  & ((Mux191) # ((Mux311 & Mux192))))

	.dataa(nRST),
	.datab(Mux31),
	.datac(Mux191),
	.datad(Mux19),
	.cin(gnd),
	.combout(\daddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~13 .lut_mask = 16'hAA80;
defparam \daddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N6
cycloneive_lcell_comb \daddr~14 (
// Equation(s):
// \daddr~14_combout  = (\nRST~input_o  & ((Mux161) # ((Mux311 & Mux162))))

	.dataa(nRST),
	.datab(Mux31),
	.datac(Mux161),
	.datad(Mux16),
	.cin(gnd),
	.combout(\daddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~14 .lut_mask = 16'hAA80;
defparam \daddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N16
cycloneive_lcell_comb \daddr~15 (
// Equation(s):
// \daddr~15_combout  = (\nRST~input_o  & ((Mux171) # ((Mux311 & Mux172))))

	.dataa(nRST),
	.datab(Mux31),
	.datac(Mux171),
	.datad(Mux17),
	.cin(gnd),
	.combout(\daddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~15 .lut_mask = 16'hAA80;
defparam \daddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N4
cycloneive_lcell_comb \daddr~16 (
// Equation(s):
// \daddr~16_combout  = (\nRST~input_o  & ((Mux141) # ((Mux311 & Mux142))))

	.dataa(nRST),
	.datab(Mux31),
	.datac(Mux14),
	.datad(Mux141),
	.cin(gnd),
	.combout(\daddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~16 .lut_mask = 16'hA8A0;
defparam \daddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N22
cycloneive_lcell_comb \daddr~17 (
// Equation(s):
// \daddr~17_combout  = (\nRST~input_o  & ((Mux151) # ((Mux311 & Mux152))))

	.dataa(Mux31),
	.datab(Mux151),
	.datac(Mux15),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~17 .lut_mask = 16'hF800;
defparam \daddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N14
cycloneive_lcell_comb \daddr~18 (
// Equation(s):
// \daddr~18_combout  = (\nRST~input_o  & ((Mux121) # ((Mux122 & Mux311))))

	.dataa(nRST),
	.datab(Mux121),
	.datac(Mux31),
	.datad(Mux12),
	.cin(gnd),
	.combout(\daddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~18 .lut_mask = 16'hAA80;
defparam \daddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N26
cycloneive_lcell_comb \daddr~19 (
// Equation(s):
// \daddr~19_combout  = (\nRST~input_o  & ((Mux131) # ((Mux311 & Mux132))))

	.dataa(nRST),
	.datab(Mux31),
	.datac(Mux131),
	.datad(Mux13),
	.cin(gnd),
	.combout(\daddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~19 .lut_mask = 16'hAA80;
defparam \daddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N16
cycloneive_lcell_comb \daddr~20 (
// Equation(s):
// \daddr~20_combout  = (\nRST~input_o  & ((Mux101) # ((Mux311 & Mux102))))

	.dataa(Mux31),
	.datab(Mux101),
	.datac(nRST),
	.datad(Mux10),
	.cin(gnd),
	.combout(\daddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~20 .lut_mask = 16'hF080;
defparam \daddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N24
cycloneive_lcell_comb \daddr~21 (
// Equation(s):
// \daddr~21_combout  = (\nRST~input_o  & ((Mux112) # ((Mux113 & Mux311))))

	.dataa(Mux112),
	.datab(Mux31),
	.datac(nRST),
	.datad(Mux111),
	.cin(gnd),
	.combout(\daddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~21 .lut_mask = 16'hF080;
defparam \daddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N20
cycloneive_lcell_comb \daddr~22 (
// Equation(s):
// \daddr~22_combout  = (\nRST~input_o  & Mux81)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Mux8),
	.cin(gnd),
	.combout(\daddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~22 .lut_mask = 16'hCC00;
defparam \daddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N10
cycloneive_lcell_comb \daddr~23 (
// Equation(s):
// \daddr~23_combout  = (\nRST~input_o  & ((Mux91) # ((Mux311 & Mux92))))

	.dataa(nRST),
	.datab(Mux31),
	.datac(Mux91),
	.datad(Mux9),
	.cin(gnd),
	.combout(\daddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~23 .lut_mask = 16'hAA80;
defparam \daddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N4
cycloneive_lcell_comb \daddr~24 (
// Equation(s):
// \daddr~24_combout  = (!Selector0 & (\nRST~input_o  & Mux64))

	.dataa(Selector0),
	.datab(nRST),
	.datac(gnd),
	.datad(Mux6),
	.cin(gnd),
	.combout(\daddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~24 .lut_mask = 16'h4400;
defparam \daddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N16
cycloneive_lcell_comb \daddr~25 (
// Equation(s):
// \daddr~25_combout  = (\nRST~input_o  & (!Selector0 & Mux71))

	.dataa(nRST),
	.datab(Selector0),
	.datac(gnd),
	.datad(Mux7),
	.cin(gnd),
	.combout(\daddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~25 .lut_mask = 16'h2200;
defparam \daddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N6
cycloneive_lcell_comb \daddr~26 (
// Equation(s):
// \daddr~26_combout  = (\nRST~input_o  & (Mux410 & !Selector0))

	.dataa(gnd),
	.datab(nRST),
	.datac(Mux4),
	.datad(Selector0),
	.cin(gnd),
	.combout(\daddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~26 .lut_mask = 16'h00C0;
defparam \daddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N2
cycloneive_lcell_comb \daddr~27 (
// Equation(s):
// \daddr~27_combout  = (\nRST~input_o  & (Mux510 & !Selector0))

	.dataa(gnd),
	.datab(nRST),
	.datac(Mux5),
	.datad(Selector0),
	.cin(gnd),
	.combout(\daddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~27 .lut_mask = 16'h00C0;
defparam \daddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N8
cycloneive_lcell_comb \daddr~28 (
// Equation(s):
// \daddr~28_combout  = (\nRST~input_o  & Mux210)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Mux2),
	.cin(gnd),
	.combout(\daddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~28 .lut_mask = 16'hF000;
defparam \daddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N30
cycloneive_lcell_comb \daddr~29 (
// Equation(s):
// \daddr~29_combout  = (\nRST~input_o  & Mux310)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Mux3),
	.cin(gnd),
	.combout(\daddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~29 .lut_mask = 16'hF000;
defparam \daddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N4
cycloneive_lcell_comb \daddr~30 (
// Equation(s):
// \daddr~30_combout  = (\nRST~input_o  & ((Mux01) # ((Mux311 & Mux02))))

	.dataa(nRST),
	.datab(Mux31),
	.datac(Mux01),
	.datad(Mux0),
	.cin(gnd),
	.combout(\daddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~30 .lut_mask = 16'hAA80;
defparam \daddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N24
cycloneive_lcell_comb \daddr~31 (
// Equation(s):
// \daddr~31_combout  = (\nRST~input_o  & ((Mux110) # ((Mux111 & Mux311))))

	.dataa(Mux11),
	.datab(Mux31),
	.datac(nRST),
	.datad(Mux1),
	.cin(gnd),
	.combout(\daddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~31 .lut_mask = 16'hF080;
defparam \daddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N14
cycloneive_lcell_comb \instr~1 (
// Equation(s):
// \instr~1_combout  = (\nRST~input_o  & (always03 & (LessThan1 & ramiframload_26)))

	.dataa(nRST),
	.datab(always0),
	.datac(LessThan1),
	.datad(ramiframload_26),
	.cin(gnd),
	.combout(\instr~1_combout ),
	.cout());
// synopsys translate_off
defparam \instr~1 .lut_mask = 16'h8000;
defparam \instr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N3
dffeas \instr[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[26] .is_wysiwyg = "true";
defparam \instr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N12
cycloneive_lcell_comb \instr~2 (
// Equation(s):
// \instr~2_combout  = (\nRST~input_o  & ((ramiframload_27) # ((!LessThan1) # (!always03))))

	.dataa(ramiframload_27),
	.datab(always0),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~2_combout ),
	.cout());
// synopsys translate_off
defparam \instr~2 .lut_mask = 16'hBF00;
defparam \instr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N29
dffeas \instr[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[27] .is_wysiwyg = "true";
defparam \instr[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N2
cycloneive_lcell_comb \instr~3 (
// Equation(s):
// \instr~3_combout  = (\nRST~input_o  & ((ramiframload_28) # ((!LessThan1) # (!always03))))

	.dataa(ramiframload_28),
	.datab(always0),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~3_combout ),
	.cout());
// synopsys translate_off
defparam \instr~3 .lut_mask = 16'hBF00;
defparam \instr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N15
dffeas \instr[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[28] .is_wysiwyg = "true";
defparam \instr[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N2
cycloneive_lcell_comb \instr~4 (
// Equation(s):
// \instr~4_combout  = (\nRST~input_o  & (((ramiframload_29) # (!LessThan1)) # (!always03)))

	.dataa(always0),
	.datab(ramiframload_29),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~4_combout ),
	.cout());
// synopsys translate_off
defparam \instr~4 .lut_mask = 16'hDF00;
defparam \instr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N9
dffeas \instr[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[29] .is_wysiwyg = "true";
defparam \instr[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N0
cycloneive_lcell_comb \instr~5 (
// Equation(s):
// \instr~5_combout  = (\nRST~input_o  & (always03 & (LessThan1 & ramiframload_30)))

	.dataa(nRST),
	.datab(always0),
	.datac(LessThan1),
	.datad(ramiframload_30),
	.cin(gnd),
	.combout(\instr~5_combout ),
	.cout());
// synopsys translate_off
defparam \instr~5 .lut_mask = 16'h8000;
defparam \instr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N19
dffeas \instr[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[30] .is_wysiwyg = "true";
defparam \instr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N24
cycloneive_lcell_comb \instr~6 (
// Equation(s):
// \instr~6_combout  = (\nRST~input_o  & (((ramiframload_31) # (!LessThan1)) # (!always03)))

	.dataa(always0),
	.datab(nRST),
	.datac(LessThan1),
	.datad(ramiframload_31),
	.cin(gnd),
	.combout(\instr~6_combout ),
	.cout());
// synopsys translate_off
defparam \instr~6 .lut_mask = 16'hCC4C;
defparam \instr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N5
dffeas \instr[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[31] .is_wysiwyg = "true";
defparam \instr[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N4
cycloneive_lcell_comb \instr~7 (
// Equation(s):
// \instr~7_combout  = (ramiframload_19 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_19),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~7_combout ),
	.cout());
// synopsys translate_off
defparam \instr~7 .lut_mask = 16'hCC00;
defparam \instr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N31
dffeas \instr[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[19] .is_wysiwyg = "true";
defparam \instr[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N16
cycloneive_lcell_comb \instr~8 (
// Equation(s):
// \instr~8_combout  = (ramiframload_18 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_18),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~8_combout ),
	.cout());
// synopsys translate_off
defparam \instr~8 .lut_mask = 16'hCC00;
defparam \instr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N27
dffeas \instr[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[18] .is_wysiwyg = "true";
defparam \instr[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N22
cycloneive_lcell_comb \instr~9 (
// Equation(s):
// \instr~9_combout  = (\nRST~input_o  & (((ramiframload_16) # (!LessThan1)) # (!always03)))

	.dataa(nRST),
	.datab(always0),
	.datac(LessThan1),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(\instr~9_combout ),
	.cout());
// synopsys translate_off
defparam \instr~9 .lut_mask = 16'hAA2A;
defparam \instr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N5
dffeas \instr[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[16] .is_wysiwyg = "true";
defparam \instr[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N18
cycloneive_lcell_comb \instr~10 (
// Equation(s):
// \instr~10_combout  = (ramiframload_17 & (\nRST~input_o  & (LessThan1 & always03)))

	.dataa(ramiframload_17),
	.datab(nRST),
	.datac(LessThan1),
	.datad(always0),
	.cin(gnd),
	.combout(\instr~10_combout ),
	.cout());
// synopsys translate_off
defparam \instr~10 .lut_mask = 16'h8000;
defparam \instr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N15
dffeas \instr[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[17] .is_wysiwyg = "true";
defparam \instr[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N30
cycloneive_lcell_comb \instr~11 (
// Equation(s):
// \instr~11_combout  = (ramiframload_20 & \nRST~input_o )

	.dataa(ramiframload_20),
	.datab(gnd),
	.datac(nRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~11_combout ),
	.cout());
// synopsys translate_off
defparam \instr~11 .lut_mask = 16'hA0A0;
defparam \instr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N13
dffeas \instr[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[20] .is_wysiwyg = "true";
defparam \instr[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N4
cycloneive_lcell_comb \instr~12 (
// Equation(s):
// \instr~12_combout  = (\nRST~input_o  & ramiframload_24)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(ramiframload_24),
	.cin(gnd),
	.combout(\instr~12_combout ),
	.cout());
// synopsys translate_off
defparam \instr~12 .lut_mask = 16'hCC00;
defparam \instr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N27
dffeas \instr[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[24] .is_wysiwyg = "true";
defparam \instr[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N10
cycloneive_lcell_comb \instr~13 (
// Equation(s):
// \instr~13_combout  = (\nRST~input_o  & ramiframload_23)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(\instr~13_combout ),
	.cout());
// synopsys translate_off
defparam \instr~13 .lut_mask = 16'hCC00;
defparam \instr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N13
dffeas \instr[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[23] .is_wysiwyg = "true";
defparam \instr[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N22
cycloneive_lcell_comb \instr~14 (
// Equation(s):
// \instr~14_combout  = (ramiframload_211 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_21),
	.datac(nRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~14_combout ),
	.cout());
// synopsys translate_off
defparam \instr~14 .lut_mask = 16'hC0C0;
defparam \instr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N5
dffeas \instr[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[21] .is_wysiwyg = "true";
defparam \instr[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N8
cycloneive_lcell_comb \instr~15 (
// Equation(s):
// \instr~15_combout  = (\nRST~input_o  & ramiframload_22)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(ramiframload_22),
	.cin(gnd),
	.combout(\instr~15_combout ),
	.cout());
// synopsys translate_off
defparam \instr~15 .lut_mask = 16'hF000;
defparam \instr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N17
dffeas \instr[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[22] .is_wysiwyg = "true";
defparam \instr[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N16
cycloneive_lcell_comb \instr~16 (
// Equation(s):
// \instr~16_combout  = (ramiframload_25 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_25),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~16_combout ),
	.cout());
// synopsys translate_off
defparam \instr~16 .lut_mask = 16'hCC00;
defparam \instr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N21
dffeas \instr[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[25] .is_wysiwyg = "true";
defparam \instr[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N30
cycloneive_lcell_comb \instr~17 (
// Equation(s):
// \instr~17_combout  = (ramiframload_3 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_3),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~17_combout ),
	.cout());
// synopsys translate_off
defparam \instr~17 .lut_mask = 16'hCC00;
defparam \instr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N31
dffeas \instr[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[3] .is_wysiwyg = "true";
defparam \instr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N10
cycloneive_lcell_comb \instr~18 (
// Equation(s):
// \instr~18_combout  = (\nRST~input_o  & (((ramiframload_4) # (!LessThan1)) # (!always03)))

	.dataa(always0),
	.datab(ramiframload_4),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~18_combout ),
	.cout());
// synopsys translate_off
defparam \instr~18 .lut_mask = 16'hDF00;
defparam \instr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N5
dffeas \instr[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[4] .is_wysiwyg = "true";
defparam \instr[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N26
cycloneive_lcell_comb \instr~19 (
// Equation(s):
// \instr~19_combout  = (LessThan1 & (always03 & (\nRST~input_o  & ramiframload_2)))

	.dataa(LessThan1),
	.datab(always0),
	.datac(nRST),
	.datad(ramiframload_2),
	.cin(gnd),
	.combout(\instr~19_combout ),
	.cout());
// synopsys translate_off
defparam \instr~19 .lut_mask = 16'h8000;
defparam \instr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N23
dffeas \instr[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[2] .is_wysiwyg = "true";
defparam \instr[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N28
cycloneive_lcell_comb \instr~20 (
// Equation(s):
// \instr~20_combout  = (\nRST~input_o  & (always03 & (LessThan1 & ramiframload_5)))

	.dataa(nRST),
	.datab(always0),
	.datac(LessThan1),
	.datad(ramiframload_5),
	.cin(gnd),
	.combout(\instr~20_combout ),
	.cout());
// synopsys translate_off
defparam \instr~20 .lut_mask = 16'h8000;
defparam \instr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N21
dffeas \instr[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[5] .is_wysiwyg = "true";
defparam \instr[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N26
cycloneive_lcell_comb \instr~21 (
// Equation(s):
// \instr~21_combout  = (\nRST~input_o  & ((ramiframload_0) # ((!LessThan1) # (!always03))))

	.dataa(ramiframload_0),
	.datab(always0),
	.datac(LessThan1),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~21_combout ),
	.cout());
// synopsys translate_off
defparam \instr~21 .lut_mask = 16'hBF00;
defparam \instr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N11
dffeas \instr[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[0] .is_wysiwyg = "true";
defparam \instr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N20
cycloneive_lcell_comb \instr~22 (
// Equation(s):
// \instr~22_combout  = (ramiframload_1 & \nRST~input_o )

	.dataa(ramiframload_1),
	.datab(gnd),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~22_combout ),
	.cout());
// synopsys translate_off
defparam \instr~22 .lut_mask = 16'hAA00;
defparam \instr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N15
dffeas \instr[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[1] .is_wysiwyg = "true";
defparam \instr[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N0
cycloneive_lcell_comb \instr~23 (
// Equation(s):
// \instr~23_combout  = (ramiframload_15 & \nRST~input_o )

	.dataa(ramiframload_15),
	.datab(gnd),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~23_combout ),
	.cout());
// synopsys translate_off
defparam \instr~23 .lut_mask = 16'hAA00;
defparam \instr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N25
dffeas \instr[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[15] .is_wysiwyg = "true";
defparam \instr[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N22
cycloneive_lcell_comb \instr~24 (
// Equation(s):
// \instr~24_combout  = (ramiframload_14 & \nRST~input_o )

	.dataa(ramiframload_14),
	.datab(nRST),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~24_combout ),
	.cout());
// synopsys translate_off
defparam \instr~24 .lut_mask = 16'h8888;
defparam \instr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N29
dffeas \instr[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[14] .is_wysiwyg = "true";
defparam \instr[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N8
cycloneive_lcell_comb \instr~25 (
// Equation(s):
// \instr~25_combout  = (ramiframload_13 & \nRST~input_o )

	.dataa(ramiframload_13),
	.datab(gnd),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~25_combout ),
	.cout());
// synopsys translate_off
defparam \instr~25 .lut_mask = 16'hAA00;
defparam \instr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N7
dffeas \instr[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[13] .is_wysiwyg = "true";
defparam \instr[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N10
cycloneive_lcell_comb \instr~26 (
// Equation(s):
// \instr~26_combout  = (ramiframload_12 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_12),
	.datac(nRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~26_combout ),
	.cout());
// synopsys translate_off
defparam \instr~26 .lut_mask = 16'hC0C0;
defparam \instr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N5
dffeas \instr[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[12] .is_wysiwyg = "true";
defparam \instr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N10
cycloneive_lcell_comb \instr~27 (
// Equation(s):
// \instr~27_combout  = (ramiframload_11 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_11),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~27_combout ),
	.cout());
// synopsys translate_off
defparam \instr~27 .lut_mask = 16'hCC00;
defparam \instr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N19
dffeas \instr[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[11] .is_wysiwyg = "true";
defparam \instr[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N22
cycloneive_lcell_comb \instr~28 (
// Equation(s):
// \instr~28_combout  = (ramiframload_10 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_10),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~28_combout ),
	.cout());
// synopsys translate_off
defparam \instr~28 .lut_mask = 16'hCC00;
defparam \instr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N9
dffeas \instr[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[10] .is_wysiwyg = "true";
defparam \instr[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N10
cycloneive_lcell_comb \instr~29 (
// Equation(s):
// \instr~29_combout  = (ramiframload_9 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_9),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~29_combout ),
	.cout());
// synopsys translate_off
defparam \instr~29 .lut_mask = 16'hCC00;
defparam \instr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N27
dffeas \instr[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[9] .is_wysiwyg = "true";
defparam \instr[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N14
cycloneive_lcell_comb \instr~30 (
// Equation(s):
// \instr~30_combout  = (ramiframload_8 & \nRST~input_o )

	.dataa(ramiframload_8),
	.datab(gnd),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~30_combout ),
	.cout());
// synopsys translate_off
defparam \instr~30 .lut_mask = 16'hAA00;
defparam \instr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N5
dffeas \instr[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[8] .is_wysiwyg = "true";
defparam \instr[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N6
cycloneive_lcell_comb \instr~31 (
// Equation(s):
// \instr~31_combout  = (ramiframload_7 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_7),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~31_combout ),
	.cout());
// synopsys translate_off
defparam \instr~31 .lut_mask = 16'hCC00;
defparam \instr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N23
dffeas \instr[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[7] .is_wysiwyg = "true";
defparam \instr[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N28
cycloneive_lcell_comb \instr~32 (
// Equation(s):
// \instr~32_combout  = (\nRST~input_o  & ramiframload_6)

	.dataa(nRST),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_6),
	.cin(gnd),
	.combout(\instr~32_combout ),
	.cout());
// synopsys translate_off
defparam \instr~32 .lut_mask = 16'hAA00;
defparam \instr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N21
dffeas \instr[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\instr[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[6] .is_wysiwyg = "true";
defparam \instr[6] .power_up = "low";
// synopsys translate_on

endmodule

module datapath (
	PC_29,
	PC_28,
	PC_31,
	PC_30,
	dpifhalt,
	PC_1,
	ruifdWEN_r,
	ruifdREN_r,
	PC_0,
	PC_3,
	PC_2,
	PC_5,
	PC_4,
	PC_7,
	PC_6,
	PC_9,
	PC_8,
	PC_11,
	PC_10,
	PC_13,
	PC_12,
	PC_15,
	PC_14,
	PC_17,
	PC_16,
	PC_19,
	PC_18,
	PC_21,
	PC_20,
	PC_23,
	PC_22,
	PC_25,
	PC_24,
	PC_27,
	PC_26,
	ramiframload_0,
	always1,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ccifiwait_0,
	ccifiwait_01,
	dcifimemload_26,
	dcifimemload_27,
	dcifimemload_28,
	dcifimemload_29,
	dcifimemload_30,
	dcifimemload_31,
	\dpif.ihit ,
	dcifimemload_19,
	dcifimemload_18,
	dcifimemload_16,
	dcifimemload_17,
	Mux63,
	Mux631,
	dcifimemload_20,
	dcifimemload_24,
	dcifimemload_23,
	dcifimemload_21,
	dcifimemload_22,
	dcifimemload_25,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_0,
	dcifimemload_1,
	Mux33,
	dcifimemload_15,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux36,
	Mux361,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux44,
	Mux441,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	Mux49,
	Mux491,
	dcifimemload_14,
	Mux50,
	Mux501,
	dcifimemload_13,
	Mux51,
	Mux511,
	dcifimemload_12,
	Mux52,
	Mux521,
	dcifimemload_11,
	Mux53,
	Mux531,
	dcifimemload_10,
	Mux54,
	Mux541,
	dcifimemload_9,
	Mux55,
	Mux551,
	dcifimemload_8,
	Mux56,
	Mux561,
	dcifimemload_7,
	Mux57,
	Mux571,
	dcifimemload_6,
	Mux58,
	Mux581,
	Mux59,
	Mux591,
	Mux60,
	Mux601,
	Mux61,
	Mux611,
	Mux62,
	Mux621,
	Mux32,
	Mux321,
	Selector0,
	Mux1,
	Mux31,
	Mux11,
	Mux0,
	Mux01,
	Mux24,
	Mux25,
	Mux26,
	Mux27,
	Mux4,
	Mux5,
	Mux6,
	Mux7,
	Mux3,
	Mux2,
	Mux23,
	Mux231,
	Mux22,
	Mux221,
	Mux21,
	Mux211,
	Mux20,
	Mux201,
	Mux19,
	Mux191,
	Mux18,
	Mux181,
	Mux17,
	Mux171,
	Mux16,
	Mux161,
	Mux29,
	Mux28,
	Mux8,
	Mux10,
	Mux101,
	Mux9,
	Mux91,
	Mux30,
	Mux15,
	Mux151,
	Mux14,
	Mux141,
	Mux13,
	Mux131,
	Mux12,
	Mux121,
	Mux111,
	Mux112,
	Mux311,
	CLK,
	nRST,
	dpifhalt1,
	devpor,
	devclrn,
	devoe);
output 	PC_29;
output 	PC_28;
output 	PC_31;
output 	PC_30;
output 	dpifhalt;
output 	PC_1;
output 	ruifdWEN_r;
output 	ruifdREN_r;
output 	PC_0;
output 	PC_3;
output 	PC_2;
output 	PC_5;
output 	PC_4;
output 	PC_7;
output 	PC_6;
output 	PC_9;
output 	PC_8;
output 	PC_11;
output 	PC_10;
output 	PC_13;
output 	PC_12;
output 	PC_15;
output 	PC_14;
output 	PC_17;
output 	PC_16;
output 	PC_19;
output 	PC_18;
output 	PC_21;
output 	PC_20;
output 	PC_23;
output 	PC_22;
output 	PC_25;
output 	PC_24;
output 	PC_27;
output 	PC_26;
input 	ramiframload_0;
input 	always1;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	ccifiwait_0;
input 	ccifiwait_01;
input 	dcifimemload_26;
input 	dcifimemload_27;
input 	dcifimemload_28;
input 	dcifimemload_29;
input 	dcifimemload_30;
input 	dcifimemload_31;
input 	\dpif.ihit ;
input 	dcifimemload_19;
input 	dcifimemload_18;
input 	dcifimemload_16;
input 	dcifimemload_17;
output 	Mux63;
output 	Mux631;
input 	dcifimemload_20;
input 	dcifimemload_24;
input 	dcifimemload_23;
input 	dcifimemload_21;
input 	dcifimemload_22;
input 	dcifimemload_25;
input 	dcifimemload_3;
input 	dcifimemload_4;
input 	dcifimemload_2;
input 	dcifimemload_5;
input 	dcifimemload_0;
input 	dcifimemload_1;
output 	Mux33;
input 	dcifimemload_15;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux36;
output 	Mux361;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux41;
output 	Mux411;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux44;
output 	Mux441;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux48;
output 	Mux481;
output 	Mux49;
output 	Mux491;
input 	dcifimemload_14;
output 	Mux50;
output 	Mux501;
input 	dcifimemload_13;
output 	Mux51;
output 	Mux511;
input 	dcifimemload_12;
output 	Mux52;
output 	Mux521;
input 	dcifimemload_11;
output 	Mux53;
output 	Mux531;
input 	dcifimemload_10;
output 	Mux54;
output 	Mux541;
input 	dcifimemload_9;
output 	Mux55;
output 	Mux551;
input 	dcifimemload_8;
output 	Mux56;
output 	Mux561;
input 	dcifimemload_7;
output 	Mux57;
output 	Mux571;
input 	dcifimemload_6;
output 	Mux58;
output 	Mux581;
output 	Mux59;
output 	Mux591;
output 	Mux60;
output 	Mux601;
output 	Mux61;
output 	Mux611;
output 	Mux62;
output 	Mux621;
output 	Mux32;
output 	Mux321;
output 	Selector0;
output 	Mux1;
output 	Mux31;
output 	Mux11;
output 	Mux0;
output 	Mux01;
output 	Mux24;
output 	Mux25;
output 	Mux26;
output 	Mux27;
output 	Mux4;
output 	Mux5;
output 	Mux6;
output 	Mux7;
output 	Mux3;
output 	Mux2;
output 	Mux23;
output 	Mux231;
output 	Mux22;
output 	Mux221;
output 	Mux21;
output 	Mux211;
output 	Mux20;
output 	Mux201;
output 	Mux19;
output 	Mux191;
output 	Mux18;
output 	Mux181;
output 	Mux17;
output 	Mux171;
output 	Mux16;
output 	Mux161;
output 	Mux29;
output 	Mux28;
output 	Mux8;
output 	Mux10;
output 	Mux101;
output 	Mux9;
output 	Mux91;
output 	Mux30;
output 	Mux15;
output 	Mux151;
output 	Mux14;
output 	Mux141;
output 	Mux13;
output 	Mux131;
output 	Mux12;
output 	Mux121;
output 	Mux111;
output 	Mux112;
output 	Mux311;
input 	CLK;
input 	nRST;
output 	dpifhalt1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add2~8_combout ;
wire \Add1~18_combout ;
wire \Add2~16_combout ;
wire \Add2~24_combout ;
wire \Add2~32_combout ;
wire \Add2~40_combout ;
wire \Add1~44_combout ;
wire \Add1~48_combout ;
wire \Add1~50_combout ;
wire \rf|Mux30~20_combout ;
wire \cu|Selector5~2_combout ;
wire \ru|nxtwen~4_combout ;
wire \cu|WideOr3~1_combout ;
wire \cu|cuif.ALUSrc[1]~5_combout ;
wire \Selector95~0_combout ;
wire \cu|Decoder1~1_combout ;
wire \Equal13~0_combout ;
wire \cu|WideOr13~0_combout ;
wire \Selector84~0_combout ;
wire \Selector95~1_combout ;
wire \Selector70~0_combout ;
wire \cu|Selector3~3_combout ;
wire \rf|Mux1~20_combout ;
wire \Selector71~0_combout ;
wire \rf|Mux2~20_combout ;
wire \Selector72~0_combout ;
wire \rf|Mux3~20_combout ;
wire \Selector73~0_combout ;
wire \rf|Mux4~20_combout ;
wire \Selector74~0_combout ;
wire \rf|Mux5~20_combout ;
wire \Selector75~0_combout ;
wire \rf|Mux6~20_combout ;
wire \Selector76~0_combout ;
wire \rf|Mux7~20_combout ;
wire \Selector77~0_combout ;
wire \rf|Mux8~20_combout ;
wire \Selector78~0_combout ;
wire \rf|Mux9~20_combout ;
wire \Selector79~0_combout ;
wire \rf|Mux10~20_combout ;
wire \Selector80~0_combout ;
wire \rf|Mux11~20_combout ;
wire \Selector81~0_combout ;
wire \rf|Mux12~20_combout ;
wire \Selector82~0_combout ;
wire \rf|Mux13~20_combout ;
wire \Selector83~0_combout ;
wire \rf|Mux14~20_combout ;
wire \Selector84~1_combout ;
wire \rf|Mux15~20_combout ;
wire \Selector85~0_combout ;
wire \rf|Mux16~20_combout ;
wire \Selector86~0_combout ;
wire \rf|Mux17~20_combout ;
wire \Selector87~0_combout ;
wire \rf|Mux18~20_combout ;
wire \Selector88~0_combout ;
wire \rf|Mux19~20_combout ;
wire \Selector89~0_combout ;
wire \rf|Mux20~20_combout ;
wire \Selector90~0_combout ;
wire \rf|Mux21~20_combout ;
wire \Selector91~0_combout ;
wire \rf|Mux22~20_combout ;
wire \Selector92~0_combout ;
wire \rf|Mux23~20_combout ;
wire \Selector93~0_combout ;
wire \rf|Mux24~20_combout ;
wire \Selector94~0_combout ;
wire \rf|Mux25~20_combout ;
wire \Selector95~2_combout ;
wire \rf|Mux26~20_combout ;
wire \Selector100~0_combout ;
wire \Selector96~0_combout ;
wire \Selector100~1_combout ;
wire \Selector96~1_combout ;
wire \rf|Mux27~20_combout ;
wire \Selector97~0_combout ;
wire \Selector97~1_combout ;
wire \rf|Mux28~20_combout ;
wire \Selector98~0_combout ;
wire \Selector98~1_combout ;
wire \rf|Mux29~20_combout ;
wire \Selector99~0_combout ;
wire \Selector99~1_combout ;
wire \Selector100~2_combout ;
wire \Selector100~3_combout ;
wire \rf|Mux31~20_combout ;
wire \Selector99~2_combout ;
wire \Selector100~4_combout ;
wire \Selector98~2_combout ;
wire \Selector95~3_combout ;
wire \Selector94~1_combout ;
wire \Selector93~1_combout ;
wire \Selector92~1_combout ;
wire \Selector91~1_combout ;
wire \Selector90~1_combout ;
wire \Selector89~1_combout ;
wire \Selector88~1_combout ;
wire \Selector87~1_combout ;
wire \Selector86~1_combout ;
wire \Selector85~1_combout ;
wire \Selector84~2_combout ;
wire \Selector83~1_combout ;
wire \Selector82~1_combout ;
wire \Selector81~1_combout ;
wire \Selector80~1_combout ;
wire \Selector79~1_combout ;
wire \Selector78~1_combout ;
wire \Selector77~1_combout ;
wire \Selector76~1_combout ;
wire \Selector75~1_combout ;
wire \Selector74~1_combout ;
wire \Selector73~1_combout ;
wire \Selector72~1_combout ;
wire \Selector71~1_combout ;
wire \Selector70~1_combout ;
wire \Selector69~0_combout ;
wire \Selector69~1_combout ;
wire \Selector96~2_combout ;
wire \rf|Mux0~20_combout ;
wire \Selector97~2_combout ;
wire \cu|Selector1~3_combout ;
wire \cu|Selector2~1_combout ;
wire \ALU|Equal0~2_combout ;
wire \ALU|Equal0~10_combout ;
wire \cu|Selector6~1_combout ;
wire \cu|cuif.RegSel[0]~3_combout ;
wire \cu|cuif.RegSel[1]~4_combout ;
wire \cu|Decoder1~2_combout ;
wire \Selector68~0_combout ;
wire \Equal10~0_combout ;
wire \Selector68~1_combout ;
wire \Selector67~0_combout ;
wire \Selector64~0_combout ;
wire \Selector66~0_combout ;
wire \Selector65~0_combout ;
wire \cu|Selector4~0_combout ;
wire \cu|Selector4~2_combout ;
wire \cu|Selector4~3_combout ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector3~0_combout ;
wire \Selector3~1_combout ;
wire \Selector8~0_combout ;
wire \Selector8~1_combout ;
wire \Selector9~0_combout ;
wire \Selector9~1_combout ;
wire \Selector10~0_combout ;
wire \Selector10~1_combout ;
wire \Selector11~0_combout ;
wire \Selector11~1_combout ;
wire \Selector12~0_combout ;
wire \Selector12~1_combout ;
wire \Selector13~0_combout ;
wire \Selector13~1_combout ;
wire \Selector14~0_combout ;
wire \Selector14~1_combout ;
wire \Selector15~0_combout ;
wire \Selector15~1_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \ALU|Mux1~9_combout ;
wire \ALU|Mux0~15_combout ;
wire \ALU|Mux23~9_combout ;
wire \ALU|Mux22~7_combout ;
wire \ALU|Mux21~7_combout ;
wire \ALU|Mux20~7_combout ;
wire \ALU|Mux19~7_combout ;
wire \ALU|Mux18~10_combout ;
wire \ALU|Mux17~7_combout ;
wire \ALU|Mux16~7_combout ;
wire \ALU|Mux10~7_combout ;
wire \ALU|Mux9~9_combout ;
wire \ALU|Mux15~8_combout ;
wire \ALU|Mux14~9_combout ;
wire \ALU|Mux13~7_combout ;
wire \ALU|Mux12~7_combout ;
wire \ALU|Mux11~7_combout ;
wire \cu|cuif.RegSel[1]~5_combout ;
wire \Add1~1 ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~54_combout ;
wire \PC[29]~1_combout ;
wire \Add1~42_combout ;
wire \Add1~40_combout ;
wire \Add1~38_combout ;
wire \Add1~36_combout ;
wire \Add1~34_combout ;
wire \Add1~32_combout ;
wire \Add1~30_combout ;
wire \Add1~26_combout ;
wire \Add1~22_combout ;
wire \Add1~20_combout ;
wire \Add1~16_combout ;
wire \Add1~14_combout ;
wire \Add1~12_combout ;
wire \Add1~10_combout ;
wire \Add1~8_combout ;
wire \Add1~6_combout ;
wire \Add1~4_combout ;
wire \Add1~0_combout ;
wire \Add2~1 ;
wire \Add2~3 ;
wire \Add2~5 ;
wire \Add2~7 ;
wire \Add2~9 ;
wire \Add2~11 ;
wire \Add2~13 ;
wire \Add2~15 ;
wire \Add2~17 ;
wire \Add2~19 ;
wire \Add2~21 ;
wire \Add2~23 ;
wire \Add2~25 ;
wire \Add2~27 ;
wire \Add2~29 ;
wire \Add2~31 ;
wire \Add2~33 ;
wire \Add2~35 ;
wire \Add2~37 ;
wire \Add2~39 ;
wire \Add2~41 ;
wire \Add2~43 ;
wire \Add2~45 ;
wire \Add2~47 ;
wire \Add2~49 ;
wire \Add2~51 ;
wire \Add2~53 ;
wire \Add2~54_combout ;
wire \PC[28]~8_combout ;
wire \Add1~52_combout ;
wire \PC[28]~0_combout ;
wire \Add2~52_combout ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~58_combout ;
wire \PC[31]~3_combout ;
wire \Add2~55 ;
wire \Add2~57 ;
wire \Add2~58_combout ;
wire \Add1~56_combout ;
wire \PC[30]~2_combout ;
wire \Add2~56_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \PC[0]~9_combout ;
wire \PC[1]~6_combout ;
wire \PC[0]~7_combout ;
wire \Add1~2_combout ;
wire \Selector60~0_combout ;
wire \Add2~2_combout ;
wire \Selector60~1_combout ;
wire \Add2~0_combout ;
wire \Selector61~0_combout ;
wire \Selector61~1_combout ;
wire \Add2~6_combout ;
wire \Selector58~0_combout ;
wire \Selector58~1_combout ;
wire \Add2~4_combout ;
wire \Selector59~0_combout ;
wire \Selector59~1_combout ;
wire \Add2~10_combout ;
wire \Selector56~0_combout ;
wire \Selector56~1_combout ;
wire \Selector57~0_combout ;
wire \Selector57~1_combout ;
wire \Add2~14_combout ;
wire \Selector54~0_combout ;
wire \Selector54~1_combout ;
wire \Add2~12_combout ;
wire \Selector55~0_combout ;
wire \Selector55~1_combout ;
wire \Add2~18_combout ;
wire \Selector52~0_combout ;
wire \Selector52~1_combout ;
wire \Selector53~0_combout ;
wire \Selector53~1_combout ;
wire \Add2~22_combout ;
wire \Selector50~0_combout ;
wire \Selector50~1_combout ;
wire \Add2~20_combout ;
wire \Selector51~0_combout ;
wire \Selector51~1_combout ;
wire \Add2~26_combout ;
wire \Selector48~0_combout ;
wire \Selector48~1_combout ;
wire \Add1~24_combout ;
wire \Selector49~0_combout ;
wire \Selector49~1_combout ;
wire \Add2~30_combout ;
wire \Selector46~0_combout ;
wire \Selector46~1_combout ;
wire \Add1~28_combout ;
wire \Add2~28_combout ;
wire \Selector47~0_combout ;
wire \Selector47~1_combout ;
wire \Add2~34_combout ;
wire \Selector44~0_combout ;
wire \Selector44~1_combout ;
wire \Selector45~0_combout ;
wire \Selector45~1_combout ;
wire \Add2~38_combout ;
wire \Selector42~0_combout ;
wire \Selector42~1_combout ;
wire \Add2~36_combout ;
wire \Selector43~0_combout ;
wire \Selector43~1_combout ;
wire \Add2~42_combout ;
wire \Selector40~0_combout ;
wire \Selector40~1_combout ;
wire \Selector41~0_combout ;
wire \Selector41~1_combout ;
wire \Add2~46_combout ;
wire \Add1~46_combout ;
wire \Selector38~0_combout ;
wire \Selector38~1_combout ;
wire \Add2~44_combout ;
wire \Selector39~0_combout ;
wire \Selector39~1_combout ;
wire \Add2~50_combout ;
wire \Selector36~0_combout ;
wire \Selector36~1_combout ;
wire \Add2~48_combout ;
wire \Selector37~0_combout ;
wire \Selector37~1_combout ;


request_unit ru(
	.dpifhalt(dpifhalt),
	.ruifdWEN_r(ruifdWEN_r),
	.ruifdREN_r(ruifdREN_r),
	.always1(always1),
	.dcifimemload_26(dcifimemload_26),
	.dcifimemload_27(dcifimemload_27),
	.dcifimemload_28(dcifimemload_28),
	.dcifimemload_29(dcifimemload_29),
	.dcifimemload_30(dcifimemload_30),
	.dcifimemload_31(dcifimemload_31),
	.nxtwen(\ru|nxtwen~4_combout ),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

control_unit cu(
	.always1(always1),
	.ccifiwait_0(ccifiwait_0),
	.dcifimemload_26(dcifimemload_26),
	.dcifimemload_27(dcifimemload_27),
	.dcifimemload_28(dcifimemload_28),
	.dcifimemload_29(dcifimemload_29),
	.dcifimemload_30(dcifimemload_30),
	.dcifimemload_31(dcifimemload_31),
	.dcifihit(\dpif.ihit ),
	.dcifimemload_3(dcifimemload_3),
	.dcifimemload_4(dcifimemload_4),
	.dcifimemload_2(dcifimemload_2),
	.dcifimemload_5(dcifimemload_5),
	.dcifimemload_0(dcifimemload_0),
	.dcifimemload_1(dcifimemload_1),
	.Selector5(\cu|Selector5~2_combout ),
	.nxtwen(\ru|nxtwen~4_combout ),
	.WideOr3(\cu|WideOr3~1_combout ),
	.cuifALUSrc_1(\cu|cuif.ALUSrc[1]~5_combout ),
	.Decoder1(\cu|Decoder1~1_combout ),
	.WideOr13(\cu|WideOr13~0_combout ),
	.Selector3(\cu|Selector3~3_combout ),
	.Selector0(Selector0),
	.Selector1(\cu|Selector1~3_combout ),
	.Selector2(\cu|Selector2~1_combout ),
	.Equal0(\ALU|Equal0~2_combout ),
	.Equal01(\ALU|Equal0~10_combout ),
	.Selector6(\cu|Selector6~1_combout ),
	.cuifRegSel_0(\cu|cuif.RegSel[0]~3_combout ),
	.cuifRegSel_1(\cu|cuif.RegSel[1]~4_combout ),
	.Decoder11(\cu|Decoder1~2_combout ),
	.Selector4(\cu|Selector4~0_combout ),
	.Selector41(\cu|Selector4~2_combout ),
	.Selector42(\cu|Selector4~3_combout ),
	.Mux1(\ALU|Mux1~9_combout ),
	.cuifRegSel_11(\cu|cuif.RegSel[1]~5_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

register_file rf(
	.Add1(\Add1~0_combout ),
	.Add11(\Add1~2_combout ),
	.Add12(\Add1~4_combout ),
	.Add13(\Add1~6_combout ),
	.Add14(\Add1~8_combout ),
	.Add15(\Add1~10_combout ),
	.Add16(\Add1~12_combout ),
	.Add17(\Add1~14_combout ),
	.Add18(\Add1~16_combout ),
	.Add19(\Add1~18_combout ),
	.Add110(\Add1~20_combout ),
	.Add111(\Add1~22_combout ),
	.Add112(\Add1~24_combout ),
	.Add113(\Add1~26_combout ),
	.Add114(\Add1~44_combout ),
	.Add115(\Add1~46_combout ),
	.Add116(\Add1~48_combout ),
	.Add117(\Add1~50_combout ),
	.PC_1(PC_1),
	.PC_0(PC_0),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.dcifimemload_30(dcifimemload_30),
	.dcifimemload_31(dcifimemload_31),
	.dcifimemload_19(dcifimemload_19),
	.dcifimemload_18(dcifimemload_18),
	.dcifimemload_16(dcifimemload_16),
	.dcifimemload_17(dcifimemload_17),
	.Mux63(Mux63),
	.Mux631(Mux631),
	.dcifimemload_24(dcifimemload_24),
	.dcifimemload_23(dcifimemload_23),
	.dcifimemload_21(dcifimemload_21),
	.dcifimemload_22(dcifimemload_22),
	.dcifimemload_25(dcifimemload_25),
	.Mux30(\rf|Mux30~20_combout ),
	.Mux33(Mux33),
	.Mux331(Mux331),
	.Mux1(\rf|Mux1~20_combout ),
	.Mux34(Mux34),
	.Mux341(Mux341),
	.Mux2(\rf|Mux2~20_combout ),
	.Mux35(Mux35),
	.Mux351(Mux351),
	.Mux3(\rf|Mux3~20_combout ),
	.Mux36(Mux36),
	.Mux361(Mux361),
	.Mux4(\rf|Mux4~20_combout ),
	.Mux37(Mux37),
	.Mux371(Mux371),
	.Mux5(\rf|Mux5~20_combout ),
	.Mux38(Mux38),
	.Mux381(Mux381),
	.Mux6(\rf|Mux6~20_combout ),
	.Mux39(Mux39),
	.Mux391(Mux391),
	.Mux7(\rf|Mux7~20_combout ),
	.Mux40(Mux40),
	.Mux401(Mux401),
	.Mux8(\rf|Mux8~20_combout ),
	.Mux41(Mux41),
	.Mux411(Mux411),
	.Mux9(\rf|Mux9~20_combout ),
	.Mux42(Mux42),
	.Mux421(Mux421),
	.Mux10(\rf|Mux10~20_combout ),
	.Mux43(Mux43),
	.Mux431(Mux431),
	.Mux11(\rf|Mux11~20_combout ),
	.Mux44(Mux44),
	.Mux441(Mux441),
	.Mux12(\rf|Mux12~20_combout ),
	.Mux45(Mux45),
	.Mux451(Mux451),
	.Mux13(\rf|Mux13~20_combout ),
	.Mux46(Mux46),
	.Mux461(Mux461),
	.Mux14(\rf|Mux14~20_combout ),
	.Mux47(Mux47),
	.Mux471(Mux471),
	.Mux15(\rf|Mux15~20_combout ),
	.Mux48(Mux48),
	.Mux481(Mux481),
	.Mux16(\rf|Mux16~20_combout ),
	.Mux49(Mux49),
	.Mux491(Mux491),
	.Mux17(\rf|Mux17~20_combout ),
	.Mux50(Mux50),
	.Mux501(Mux501),
	.Mux18(\rf|Mux18~20_combout ),
	.Mux51(Mux51),
	.Mux511(Mux511),
	.Mux19(\rf|Mux19~20_combout ),
	.Mux52(Mux52),
	.Mux521(Mux521),
	.dcifimemload_11(dcifimemload_11),
	.Mux20(\rf|Mux20~20_combout ),
	.Mux53(Mux53),
	.Mux531(Mux531),
	.dcifimemload_10(dcifimemload_10),
	.Mux21(\rf|Mux21~20_combout ),
	.Mux54(Mux54),
	.Mux541(Mux541),
	.dcifimemload_9(dcifimemload_9),
	.Mux22(\rf|Mux22~20_combout ),
	.Mux55(Mux55),
	.Mux551(Mux551),
	.dcifimemload_8(dcifimemload_8),
	.Mux23(\rf|Mux23~20_combout ),
	.Mux56(Mux56),
	.Mux561(Mux561),
	.Mux24(\rf|Mux24~20_combout ),
	.Mux57(Mux57),
	.Mux571(Mux571),
	.Mux25(\rf|Mux25~20_combout ),
	.Mux58(Mux58),
	.Mux581(Mux581),
	.Mux26(\rf|Mux26~20_combout ),
	.Mux59(Mux59),
	.Mux591(Mux591),
	.Mux27(\rf|Mux27~20_combout ),
	.Mux60(Mux60),
	.Mux601(Mux601),
	.Mux28(\rf|Mux28~20_combout ),
	.Mux61(Mux61),
	.Mux611(Mux611),
	.Mux29(\rf|Mux29~20_combout ),
	.Mux62(Mux62),
	.Mux621(Mux621),
	.Mux31(\rf|Mux31~20_combout ),
	.Mux32(Mux32),
	.Mux321(Mux321),
	.Mux0(\rf|Mux0~20_combout ),
	.Selector0(Selector0),
	.Mux241(Mux24),
	.Mux251(Mux25),
	.Mux261(Mux26),
	.Mux271(Mux27),
	.Mux410(Mux4),
	.Mux510(Mux5),
	.Mux64(Mux6),
	.Mux71(Mux7),
	.Mux291(Mux29),
	.Mux281(Mux28),
	.Mux301(Mux30),
	.Mux311(Mux311),
	.cuifRegSel_0(\cu|cuif.RegSel[0]~3_combout ),
	.cuifRegSel_1(\cu|cuif.RegSel[1]~4_combout ),
	.Selector68(\Selector68~1_combout ),
	.Selector67(\Selector67~0_combout ),
	.Selector64(\Selector64~0_combout ),
	.Selector66(\Selector66~0_combout ),
	.Selector65(\Selector65~0_combout ),
	.Selector4(\cu|Selector4~0_combout ),
	.Selector41(\cu|Selector4~2_combout ),
	.Selector42(\cu|Selector4~3_combout ),
	.Selector1(\Selector1~1_combout ),
	.Selector2(\Selector2~1_combout ),
	.Selector3(\Selector3~1_combout ),
	.Selector8(\Selector8~1_combout ),
	.Selector9(\Selector9~1_combout ),
	.Selector10(\Selector10~1_combout ),
	.Selector11(\Selector11~1_combout ),
	.Selector12(\Selector12~1_combout ),
	.Selector13(\Selector13~1_combout ),
	.Selector14(\Selector14~1_combout ),
	.Selector15(\Selector15~1_combout ),
	.Selector01(\Selector0~1_combout ),
	.Mux231(\ALU|Mux23~9_combout ),
	.Mux221(\ALU|Mux22~7_combout ),
	.Mux211(\ALU|Mux21~7_combout ),
	.Mux201(\ALU|Mux20~7_combout ),
	.Mux191(\ALU|Mux19~7_combout ),
	.Mux181(\ALU|Mux18~10_combout ),
	.Mux171(\ALU|Mux17~7_combout ),
	.Mux161(\ALU|Mux16~7_combout ),
	.cuifRegSel_11(\cu|cuif.RegSel[1]~5_combout ),
	.CLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu ALU(
	.Mux63(Mux63),
	.Mux30(\rf|Mux30~20_combout ),
	.Selector95(\Selector95~0_combout ),
	.Mux33(Mux33),
	.Selector70(\Selector70~0_combout ),
	.Selector3(\cu|Selector3~3_combout ),
	.Mux1(\rf|Mux1~20_combout ),
	.Mux34(Mux34),
	.Selector71(\Selector71~0_combout ),
	.Mux2(\rf|Mux2~20_combout ),
	.Mux35(Mux35),
	.Selector72(\Selector72~0_combout ),
	.Mux3(\rf|Mux3~20_combout ),
	.Mux36(Mux36),
	.Selector73(\Selector73~0_combout ),
	.Mux4(\rf|Mux4~20_combout ),
	.Mux37(Mux37),
	.Selector74(\Selector74~0_combout ),
	.Mux5(\rf|Mux5~20_combout ),
	.Mux38(Mux38),
	.Selector75(\Selector75~0_combout ),
	.Mux6(\rf|Mux6~20_combout ),
	.Mux39(Mux39),
	.Selector76(\Selector76~0_combout ),
	.Mux7(\rf|Mux7~20_combout ),
	.Mux40(Mux40),
	.Selector77(\Selector77~0_combout ),
	.Mux8(\rf|Mux8~20_combout ),
	.Mux41(Mux41),
	.Selector78(\Selector78~0_combout ),
	.Mux9(\rf|Mux9~20_combout ),
	.Mux42(Mux42),
	.Selector79(\Selector79~0_combout ),
	.Mux10(\rf|Mux10~20_combout ),
	.Mux43(Mux43),
	.Selector80(\Selector80~0_combout ),
	.Mux11(\rf|Mux11~20_combout ),
	.Mux44(Mux44),
	.Selector81(\Selector81~0_combout ),
	.Mux12(\rf|Mux12~20_combout ),
	.Mux45(Mux45),
	.Selector82(\Selector82~0_combout ),
	.Mux13(\rf|Mux13~20_combout ),
	.Mux46(Mux46),
	.Selector83(\Selector83~0_combout ),
	.Mux14(\rf|Mux14~20_combout ),
	.Mux47(Mux47),
	.Selector84(\Selector84~1_combout ),
	.Mux15(\rf|Mux15~20_combout ),
	.Mux48(Mux48),
	.Selector85(\Selector85~0_combout ),
	.Mux16(\rf|Mux16~20_combout ),
	.Mux49(Mux49),
	.Selector86(\Selector86~0_combout ),
	.Mux17(\rf|Mux17~20_combout ),
	.Mux50(Mux50),
	.Selector87(\Selector87~0_combout ),
	.Mux18(\rf|Mux18~20_combout ),
	.Mux51(Mux51),
	.Selector88(\Selector88~0_combout ),
	.Mux19(\rf|Mux19~20_combout ),
	.Mux52(Mux52),
	.Selector89(\Selector89~0_combout ),
	.Mux20(\rf|Mux20~20_combout ),
	.Mux53(Mux53),
	.Selector90(\Selector90~0_combout ),
	.Mux21(\rf|Mux21~20_combout ),
	.Mux54(Mux54),
	.Selector91(\Selector91~0_combout ),
	.Mux22(\rf|Mux22~20_combout ),
	.Mux55(Mux55),
	.Selector92(\Selector92~0_combout ),
	.Mux23(\rf|Mux23~20_combout ),
	.Mux56(Mux56),
	.Selector93(\Selector93~0_combout ),
	.Mux24(\rf|Mux24~20_combout ),
	.Mux57(Mux57),
	.Selector94(\Selector94~0_combout ),
	.Mux25(\rf|Mux25~20_combout ),
	.Mux58(Mux58),
	.Selector951(\Selector95~2_combout ),
	.Mux26(\rf|Mux26~20_combout ),
	.Selector100(\Selector100~0_combout ),
	.Mux59(Mux59),
	.Selector96(\Selector96~1_combout ),
	.Mux27(\rf|Mux27~20_combout ),
	.Mux60(Mux60),
	.Selector97(\Selector97~1_combout ),
	.Mux28(\rf|Mux28~20_combout ),
	.Mux61(Mux61),
	.Selector98(\Selector98~1_combout ),
	.Mux29(\rf|Mux29~20_combout ),
	.Mux62(Mux62),
	.Selector99(\Selector99~1_combout ),
	.Selector1001(\Selector100~3_combout ),
	.Mux31(\rf|Mux31~20_combout ),
	.Selector991(\Selector99~2_combout ),
	.Selector1002(\Selector100~4_combout ),
	.Selector981(\Selector98~2_combout ),
	.Selector952(\Selector95~3_combout ),
	.Selector941(\Selector94~1_combout ),
	.Selector931(\Selector93~1_combout ),
	.Selector921(\Selector92~1_combout ),
	.Selector911(\Selector91~1_combout ),
	.Selector901(\Selector90~1_combout ),
	.Selector891(\Selector89~1_combout ),
	.Selector881(\Selector88~1_combout ),
	.Selector871(\Selector87~1_combout ),
	.Selector861(\Selector86~1_combout ),
	.Selector851(\Selector85~1_combout ),
	.Selector841(\Selector84~2_combout ),
	.Selector831(\Selector83~1_combout ),
	.Selector821(\Selector82~1_combout ),
	.Selector811(\Selector81~1_combout ),
	.Selector801(\Selector80~1_combout ),
	.Selector791(\Selector79~1_combout ),
	.Selector781(\Selector78~1_combout ),
	.Selector771(\Selector77~1_combout ),
	.Selector761(\Selector76~1_combout ),
	.Selector751(\Selector75~1_combout ),
	.Selector741(\Selector74~1_combout ),
	.Selector731(\Selector73~1_combout ),
	.Selector721(\Selector72~1_combout ),
	.Selector711(\Selector71~1_combout ),
	.Selector701(\Selector70~1_combout ),
	.Selector69(\Selector69~0_combout ),
	.Mux32(Mux321),
	.Selector691(\Selector69~1_combout ),
	.Selector961(\Selector96~2_combout ),
	.Mux0(\rf|Mux0~20_combout ),
	.Selector971(\Selector97~2_combout ),
	.Selector0(Selector0),
	.Selector1(\cu|Selector1~3_combout ),
	.Selector2(\cu|Selector2~1_combout ),
	.Mux110(Mux1),
	.Mux311(Mux31),
	.Mux111(Mux11),
	.Mux01(Mux0),
	.Mux02(Mux01),
	.Mux241(Mux24),
	.Mux251(Mux25),
	.Mux261(Mux26),
	.Mux271(Mux27),
	.Mux410(Mux4),
	.Mux510(Mux5),
	.Mux64(Mux6),
	.Mux71(Mux7),
	.Equal0(\ALU|Equal0~2_combout ),
	.Mux310(Mux3),
	.Mux210(Mux2),
	.Mux231(Mux23),
	.Mux232(Mux231),
	.Mux221(Mux22),
	.Mux222(Mux221),
	.Mux211(Mux21),
	.Mux212(Mux211),
	.Mux201(Mux20),
	.Mux202(Mux201),
	.Mux191(Mux19),
	.Mux192(Mux191),
	.Mux181(Mux18),
	.Mux182(Mux181),
	.Mux171(Mux17),
	.Mux172(Mux171),
	.Mux161(Mux16),
	.Mux162(Mux161),
	.Mux291(Mux29),
	.Mux281(Mux28),
	.Mux81(Mux8),
	.Mux101(Mux10),
	.Mux102(Mux101),
	.Mux91(Mux9),
	.Mux92(Mux91),
	.Mux301(Mux30),
	.Mux151(Mux15),
	.Mux152(Mux151),
	.Mux141(Mux14),
	.Mux142(Mux141),
	.Mux131(Mux13),
	.Mux132(Mux131),
	.Mux121(Mux12),
	.Mux122(Mux121),
	.Mux112(Mux111),
	.Mux113(Mux112),
	.Equal01(\ALU|Equal0~10_combout ),
	.Mux312(Mux311),
	.Mux114(\ALU|Mux1~9_combout ),
	.Mux03(\ALU|Mux0~15_combout ),
	.Mux233(\ALU|Mux23~9_combout ),
	.Mux223(\ALU|Mux22~7_combout ),
	.Mux213(\ALU|Mux21~7_combout ),
	.Mux203(\ALU|Mux20~7_combout ),
	.Mux193(\ALU|Mux19~7_combout ),
	.Mux183(\ALU|Mux18~10_combout ),
	.Mux173(\ALU|Mux17~7_combout ),
	.Mux163(\ALU|Mux16~7_combout ),
	.Mux103(\ALU|Mux10~7_combout ),
	.Mux93(\ALU|Mux9~9_combout ),
	.Mux153(\ALU|Mux15~8_combout ),
	.Mux143(\ALU|Mux14~9_combout ),
	.Mux133(\ALU|Mux13~7_combout ),
	.Mux123(\ALU|Mux12~7_combout ),
	.Mux115(\ALU|Mux11~7_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X66_Y42_N10
cycloneive_lcell_comb \Add2~8 (
// Equation(s):
// \Add2~8_combout  = ((dcifimemload_4 $ (\Add1~8_combout  $ (!\Add2~7 )))) # (GND)
// \Add2~9  = CARRY((dcifimemload_4 & ((\Add1~8_combout ) # (!\Add2~7 ))) # (!dcifimemload_4 & (\Add1~8_combout  & !\Add2~7 )))

	.dataa(dcifimemload_4),
	.datab(\Add1~8_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout(\Add2~9 ));
// synopsys translate_off
defparam \Add2~8 .lut_mask = 16'h698E;
defparam \Add2~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N20
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (PC_11 & (!\Add1~17 )) # (!PC_11 & ((\Add1~17 ) # (GND)))
// \Add1~19  = CARRY((!\Add1~17 ) # (!PC_11))

	.dataa(PC_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h5A5F;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N18
cycloneive_lcell_comb \Add2~16 (
// Equation(s):
// \Add2~16_combout  = ((dcifimemload_8 $ (\Add1~16_combout  $ (!\Add2~15 )))) # (GND)
// \Add2~17  = CARRY((dcifimemload_8 & ((\Add1~16_combout ) # (!\Add2~15 ))) # (!dcifimemload_8 & (\Add1~16_combout  & !\Add2~15 )))

	.dataa(dcifimemload_8),
	.datab(\Add1~16_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~15 ),
	.combout(\Add2~16_combout ),
	.cout(\Add2~17 ));
// synopsys translate_off
defparam \Add2~16 .lut_mask = 16'h698E;
defparam \Add2~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N26
cycloneive_lcell_comb \Add2~24 (
// Equation(s):
// \Add2~24_combout  = ((\Add1~24_combout  $ (dcifimemload_12 $ (!\Add2~23 )))) # (GND)
// \Add2~25  = CARRY((\Add1~24_combout  & ((dcifimemload_12) # (!\Add2~23 ))) # (!\Add1~24_combout  & (dcifimemload_12 & !\Add2~23 )))

	.dataa(\Add1~24_combout ),
	.datab(dcifimemload_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~23 ),
	.combout(\Add2~24_combout ),
	.cout(\Add2~25 ));
// synopsys translate_off
defparam \Add2~24 .lut_mask = 16'h698E;
defparam \Add2~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N2
cycloneive_lcell_comb \Add2~32 (
// Equation(s):
// \Add2~32_combout  = ((dcifimemload_15 $ (\Add1~32_combout  $ (!\Add2~31 )))) # (GND)
// \Add2~33  = CARRY((dcifimemload_15 & ((\Add1~32_combout ) # (!\Add2~31 ))) # (!dcifimemload_15 & (\Add1~32_combout  & !\Add2~31 )))

	.dataa(dcifimemload_15),
	.datab(\Add1~32_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~31 ),
	.combout(\Add2~32_combout ),
	.cout(\Add2~33 ));
// synopsys translate_off
defparam \Add2~32 .lut_mask = 16'h698E;
defparam \Add2~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N10
cycloneive_lcell_comb \Add2~40 (
// Equation(s):
// \Add2~40_combout  = ((dcifimemload_15 $ (\Add1~40_combout  $ (!\Add2~39 )))) # (GND)
// \Add2~41  = CARRY((dcifimemload_15 & ((\Add1~40_combout ) # (!\Add2~39 ))) # (!dcifimemload_15 & (\Add1~40_combout  & !\Add2~39 )))

	.dataa(dcifimemload_15),
	.datab(\Add1~40_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~39 ),
	.combout(\Add2~40_combout ),
	.cout(\Add2~41 ));
// synopsys translate_off
defparam \Add2~40 .lut_mask = 16'h698E;
defparam \Add2~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N14
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = (PC_24 & (\Add1~43  $ (GND))) # (!PC_24 & (!\Add1~43  & VCC))
// \Add1~45  = CARRY((PC_24 & !\Add1~43 ))

	.dataa(gnd),
	.datab(PC_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'hC30C;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N18
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = (PC_26 & (\Add1~47  $ (GND))) # (!PC_26 & (!\Add1~47  & VCC))
// \Add1~49  = CARRY((PC_26 & !\Add1~47 ))

	.dataa(PC_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'hA50A;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N20
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (PC_27 & (!\Add1~49 )) # (!PC_27 & ((\Add1~49 ) # (GND)))
// \Add1~51  = CARRY((!\Add1~49 ) # (!PC_27))

	.dataa(gnd),
	.datab(PC_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h3C3F;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N28
cycloneive_lcell_comb \Selector95~0 (
// Equation(s):
// \Selector95~0_combout  = (!WideOr3 & (dcifimemload_20 & !cuifALUSrc_1))

	.dataa(gnd),
	.datab(\cu|WideOr3~1_combout ),
	.datac(dcifimemload_20),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector95~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector95~0 .lut_mask = 16'h0030;
defparam \Selector95~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N18
cycloneive_lcell_comb \Equal13~0 (
// Equation(s):
// \Equal13~0_combout  = (WideOr3 & !cuifALUSrc_1)

	.dataa(gnd),
	.datab(gnd),
	.datac(\cu|WideOr3~1_combout ),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Equal13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal13~0 .lut_mask = 16'h00F0;
defparam \Equal13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N0
cycloneive_lcell_comb \Selector84~0 (
// Equation(s):
// \Selector84~0_combout  = (WideOr13 & (dcifimemload_15 & (Decoder1 & \Equal13~0_combout )))

	.dataa(\cu|WideOr13~0_combout ),
	.datab(dcifimemload_15),
	.datac(\cu|Decoder1~1_combout ),
	.datad(\Equal13~0_combout ),
	.cin(gnd),
	.combout(\Selector84~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector84~0 .lut_mask = 16'h8000;
defparam \Selector84~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N4
cycloneive_lcell_comb \Selector95~1 (
// Equation(s):
// \Selector95~1_combout  = (!dcifimemload_20 & (!WideOr3 & !cuifALUSrc_1))

	.dataa(dcifimemload_20),
	.datab(\cu|WideOr3~1_combout ),
	.datac(gnd),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector95~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector95~1 .lut_mask = 16'h0011;
defparam \Selector95~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N16
cycloneive_lcell_comb \Selector70~0 (
// Equation(s):
// \Selector70~0_combout  = (\Selector84~0_combout ) # ((\Selector95~1_combout  & Mux331))

	.dataa(gnd),
	.datab(\Selector95~1_combout ),
	.datac(Mux331),
	.datad(\Selector84~0_combout ),
	.cin(gnd),
	.combout(\Selector70~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector70~0 .lut_mask = 16'hFFC0;
defparam \Selector70~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N14
cycloneive_lcell_comb \Selector71~0 (
// Equation(s):
// \Selector71~0_combout  = (\Selector84~0_combout ) # ((Mux341 & \Selector95~1_combout ))

	.dataa(gnd),
	.datab(Mux341),
	.datac(\Selector95~1_combout ),
	.datad(\Selector84~0_combout ),
	.cin(gnd),
	.combout(\Selector71~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector71~0 .lut_mask = 16'hFFC0;
defparam \Selector71~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N0
cycloneive_lcell_comb \Selector72~0 (
// Equation(s):
// \Selector72~0_combout  = (\Selector84~0_combout ) # ((\Selector95~1_combout  & Mux351))

	.dataa(gnd),
	.datab(\Selector95~1_combout ),
	.datac(\Selector84~0_combout ),
	.datad(Mux351),
	.cin(gnd),
	.combout(\Selector72~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector72~0 .lut_mask = 16'hFCF0;
defparam \Selector72~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N14
cycloneive_lcell_comb \Selector73~0 (
// Equation(s):
// \Selector73~0_combout  = (\Selector84~0_combout ) # ((Mux361 & \Selector95~1_combout ))

	.dataa(Mux361),
	.datab(gnd),
	.datac(\Selector95~1_combout ),
	.datad(\Selector84~0_combout ),
	.cin(gnd),
	.combout(\Selector73~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector73~0 .lut_mask = 16'hFFA0;
defparam \Selector73~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N2
cycloneive_lcell_comb \Selector74~0 (
// Equation(s):
// \Selector74~0_combout  = (\Selector84~0_combout ) # ((\Selector95~1_combout  & Mux371))

	.dataa(\Selector95~1_combout ),
	.datab(gnd),
	.datac(Mux371),
	.datad(\Selector84~0_combout ),
	.cin(gnd),
	.combout(\Selector74~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector74~0 .lut_mask = 16'hFFA0;
defparam \Selector74~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N8
cycloneive_lcell_comb \Selector75~0 (
// Equation(s):
// \Selector75~0_combout  = (\Selector84~0_combout ) # ((Mux381 & \Selector95~1_combout ))

	.dataa(Mux381),
	.datab(\Selector84~0_combout ),
	.datac(gnd),
	.datad(\Selector95~1_combout ),
	.cin(gnd),
	.combout(\Selector75~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector75~0 .lut_mask = 16'hEECC;
defparam \Selector75~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N8
cycloneive_lcell_comb \Selector76~0 (
// Equation(s):
// \Selector76~0_combout  = (\Selector84~0_combout ) # ((Mux391 & \Selector95~1_combout ))

	.dataa(Mux391),
	.datab(gnd),
	.datac(\Selector95~1_combout ),
	.datad(\Selector84~0_combout ),
	.cin(gnd),
	.combout(\Selector76~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector76~0 .lut_mask = 16'hFFA0;
defparam \Selector76~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N14
cycloneive_lcell_comb \Selector77~0 (
// Equation(s):
// \Selector77~0_combout  = (\Selector84~0_combout ) # ((\Selector95~1_combout  & Mux401))

	.dataa(\Selector84~0_combout ),
	.datab(gnd),
	.datac(\Selector95~1_combout ),
	.datad(Mux401),
	.cin(gnd),
	.combout(\Selector77~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector77~0 .lut_mask = 16'hFAAA;
defparam \Selector77~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N4
cycloneive_lcell_comb \Selector78~0 (
// Equation(s):
// \Selector78~0_combout  = (\Selector84~0_combout ) # ((\Selector95~1_combout  & Mux411))

	.dataa(\Selector84~0_combout ),
	.datab(gnd),
	.datac(\Selector95~1_combout ),
	.datad(Mux411),
	.cin(gnd),
	.combout(\Selector78~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector78~0 .lut_mask = 16'hFAAA;
defparam \Selector78~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N2
cycloneive_lcell_comb \Selector79~0 (
// Equation(s):
// \Selector79~0_combout  = (\Selector84~0_combout ) # ((Mux421 & \Selector95~1_combout ))

	.dataa(\Selector84~0_combout ),
	.datab(gnd),
	.datac(Mux421),
	.datad(\Selector95~1_combout ),
	.cin(gnd),
	.combout(\Selector79~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector79~0 .lut_mask = 16'hFAAA;
defparam \Selector79~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N14
cycloneive_lcell_comb \Selector80~0 (
// Equation(s):
// \Selector80~0_combout  = (\Selector84~0_combout ) # ((\Selector95~1_combout  & Mux431))

	.dataa(gnd),
	.datab(\Selector95~1_combout ),
	.datac(\Selector84~0_combout ),
	.datad(Mux431),
	.cin(gnd),
	.combout(\Selector80~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector80~0 .lut_mask = 16'hFCF0;
defparam \Selector80~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N20
cycloneive_lcell_comb \Selector81~0 (
// Equation(s):
// \Selector81~0_combout  = (\Selector84~0_combout ) # ((\Selector95~1_combout  & Mux441))

	.dataa(\Selector95~1_combout ),
	.datab(\Selector84~0_combout ),
	.datac(gnd),
	.datad(Mux441),
	.cin(gnd),
	.combout(\Selector81~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector81~0 .lut_mask = 16'hEECC;
defparam \Selector81~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N18
cycloneive_lcell_comb \Selector82~0 (
// Equation(s):
// \Selector82~0_combout  = (\Selector84~0_combout ) # ((\Selector95~1_combout  & Mux451))

	.dataa(\Selector95~1_combout ),
	.datab(\Selector84~0_combout ),
	.datac(gnd),
	.datad(Mux451),
	.cin(gnd),
	.combout(\Selector82~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector82~0 .lut_mask = 16'hEECC;
defparam \Selector82~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N16
cycloneive_lcell_comb \Selector83~0 (
// Equation(s):
// \Selector83~0_combout  = (\Selector84~0_combout ) # ((\Selector95~1_combout  & Mux461))

	.dataa(\Selector95~1_combout ),
	.datab(\Selector84~0_combout ),
	.datac(gnd),
	.datad(Mux461),
	.cin(gnd),
	.combout(\Selector83~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector83~0 .lut_mask = 16'hEECC;
defparam \Selector83~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N8
cycloneive_lcell_comb \Selector84~1 (
// Equation(s):
// \Selector84~1_combout  = (\Selector84~0_combout ) # ((Mux471 & \Selector95~1_combout ))

	.dataa(Mux471),
	.datab(gnd),
	.datac(\Selector84~0_combout ),
	.datad(\Selector95~1_combout ),
	.cin(gnd),
	.combout(\Selector84~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector84~1 .lut_mask = 16'hFAF0;
defparam \Selector84~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N30
cycloneive_lcell_comb \Selector85~0 (
// Equation(s):
// \Selector85~0_combout  = (dcifimemload_15 & ((\Equal13~0_combout ) # ((Mux481 & \Selector95~1_combout )))) # (!dcifimemload_15 & (Mux481 & (\Selector95~1_combout )))

	.dataa(dcifimemload_15),
	.datab(Mux481),
	.datac(\Selector95~1_combout ),
	.datad(\Equal13~0_combout ),
	.cin(gnd),
	.combout(\Selector85~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector85~0 .lut_mask = 16'hEAC0;
defparam \Selector85~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N26
cycloneive_lcell_comb \Selector86~0 (
// Equation(s):
// \Selector86~0_combout  = (dcifimemload_14 & ((\Equal13~0_combout ) # ((Mux491 & \Selector95~1_combout )))) # (!dcifimemload_14 & (((Mux491 & \Selector95~1_combout ))))

	.dataa(dcifimemload_14),
	.datab(\Equal13~0_combout ),
	.datac(Mux491),
	.datad(\Selector95~1_combout ),
	.cin(gnd),
	.combout(\Selector86~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector86~0 .lut_mask = 16'hF888;
defparam \Selector86~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N2
cycloneive_lcell_comb \Selector87~0 (
// Equation(s):
// \Selector87~0_combout  = (\Equal13~0_combout  & ((dcifimemload_13) # ((Mux501 & \Selector95~1_combout )))) # (!\Equal13~0_combout  & (((Mux501 & \Selector95~1_combout ))))

	.dataa(\Equal13~0_combout ),
	.datab(dcifimemload_13),
	.datac(Mux501),
	.datad(\Selector95~1_combout ),
	.cin(gnd),
	.combout(\Selector87~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector87~0 .lut_mask = 16'hF888;
defparam \Selector87~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N6
cycloneive_lcell_comb \Selector88~0 (
// Equation(s):
// \Selector88~0_combout  = (dcifimemload_12 & ((\Equal13~0_combout ) # ((Mux511 & \Selector95~1_combout )))) # (!dcifimemload_12 & (Mux511 & (\Selector95~1_combout )))

	.dataa(dcifimemload_12),
	.datab(Mux511),
	.datac(\Selector95~1_combout ),
	.datad(\Equal13~0_combout ),
	.cin(gnd),
	.combout(\Selector88~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector88~0 .lut_mask = 16'hEAC0;
defparam \Selector88~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N4
cycloneive_lcell_comb \Selector89~0 (
// Equation(s):
// \Selector89~0_combout  = (dcifimemload_11 & ((\Equal13~0_combout ) # ((Mux521 & \Selector95~1_combout )))) # (!dcifimemload_11 & (Mux521 & (\Selector95~1_combout )))

	.dataa(dcifimemload_11),
	.datab(Mux521),
	.datac(\Selector95~1_combout ),
	.datad(\Equal13~0_combout ),
	.cin(gnd),
	.combout(\Selector89~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector89~0 .lut_mask = 16'hEAC0;
defparam \Selector89~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N30
cycloneive_lcell_comb \Selector90~0 (
// Equation(s):
// \Selector90~0_combout  = (dcifimemload_10 & ((\Equal13~0_combout ) # ((\Selector95~1_combout  & Mux531)))) # (!dcifimemload_10 & (\Selector95~1_combout  & (Mux531)))

	.dataa(dcifimemload_10),
	.datab(\Selector95~1_combout ),
	.datac(Mux531),
	.datad(\Equal13~0_combout ),
	.cin(gnd),
	.combout(\Selector90~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector90~0 .lut_mask = 16'hEAC0;
defparam \Selector90~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N28
cycloneive_lcell_comb \Selector91~0 (
// Equation(s):
// \Selector91~0_combout  = (dcifimemload_9 & ((\Equal13~0_combout ) # ((\Selector95~1_combout  & Mux541)))) # (!dcifimemload_9 & (((\Selector95~1_combout  & Mux541))))

	.dataa(dcifimemload_9),
	.datab(\Equal13~0_combout ),
	.datac(\Selector95~1_combout ),
	.datad(Mux541),
	.cin(gnd),
	.combout(\Selector91~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector91~0 .lut_mask = 16'hF888;
defparam \Selector91~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N2
cycloneive_lcell_comb \Selector92~0 (
// Equation(s):
// \Selector92~0_combout  = (\Equal13~0_combout  & ((dcifimemload_8) # ((\Selector95~1_combout  & Mux551)))) # (!\Equal13~0_combout  & (((\Selector95~1_combout  & Mux551))))

	.dataa(\Equal13~0_combout ),
	.datab(dcifimemload_8),
	.datac(\Selector95~1_combout ),
	.datad(Mux551),
	.cin(gnd),
	.combout(\Selector92~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector92~0 .lut_mask = 16'hF888;
defparam \Selector92~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N0
cycloneive_lcell_comb \Selector93~0 (
// Equation(s):
// \Selector93~0_combout  = (dcifimemload_7 & ((\Equal13~0_combout ) # ((\Selector95~1_combout  & Mux561)))) # (!dcifimemload_7 & (\Selector95~1_combout  & ((Mux561))))

	.dataa(dcifimemload_7),
	.datab(\Selector95~1_combout ),
	.datac(\Equal13~0_combout ),
	.datad(Mux561),
	.cin(gnd),
	.combout(\Selector93~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector93~0 .lut_mask = 16'hECA0;
defparam \Selector93~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N14
cycloneive_lcell_comb \Selector94~0 (
// Equation(s):
// \Selector94~0_combout  = (dcifimemload_6 & ((\Equal13~0_combout ) # ((\Selector95~1_combout  & Mux571)))) # (!dcifimemload_6 & (\Selector95~1_combout  & ((Mux571))))

	.dataa(dcifimemload_6),
	.datab(\Selector95~1_combout ),
	.datac(\Equal13~0_combout ),
	.datad(Mux571),
	.cin(gnd),
	.combout(\Selector94~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector94~0 .lut_mask = 16'hECA0;
defparam \Selector94~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N28
cycloneive_lcell_comb \Selector95~2 (
// Equation(s):
// \Selector95~2_combout  = (WideOr3 & ((dcifimemload_5) # ((\Selector95~1_combout  & Mux581)))) # (!WideOr3 & (((\Selector95~1_combout  & Mux581))))

	.dataa(\cu|WideOr3~1_combout ),
	.datab(dcifimemload_5),
	.datac(\Selector95~1_combout ),
	.datad(Mux581),
	.cin(gnd),
	.combout(\Selector95~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector95~2 .lut_mask = 16'hF888;
defparam \Selector95~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N20
cycloneive_lcell_comb \Selector100~0 (
// Equation(s):
// \Selector100~0_combout  = (dcifimemload_20 & (WideOr3 $ (!cuifALUSrc_1)))

	.dataa(gnd),
	.datab(\cu|WideOr3~1_combout ),
	.datac(dcifimemload_20),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector100~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector100~0 .lut_mask = 16'hC030;
defparam \Selector100~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N12
cycloneive_lcell_comb \Selector96~0 (
// Equation(s):
// \Selector96~0_combout  = (WideOr3 & (dcifimemload_4 & ((!cuifALUSrc_1)))) # (!WideOr3 & (((dcifimemload_10 & cuifALUSrc_1))))

	.dataa(dcifimemload_4),
	.datab(dcifimemload_10),
	.datac(\cu|WideOr3~1_combout ),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector96~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector96~0 .lut_mask = 16'h0CA0;
defparam \Selector96~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N22
cycloneive_lcell_comb \Selector100~1 (
// Equation(s):
// \Selector100~1_combout  = WideOr3 $ (cuifALUSrc_1)

	.dataa(gnd),
	.datab(gnd),
	.datac(\cu|WideOr3~1_combout ),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector100~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector100~1 .lut_mask = 16'h0FF0;
defparam \Selector100~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N28
cycloneive_lcell_comb \Selector96~1 (
// Equation(s):
// \Selector96~1_combout  = (\Selector96~0_combout ) # ((Mux591 & (!dcifimemload_20 & !\Selector100~1_combout )))

	.dataa(\Selector96~0_combout ),
	.datab(Mux591),
	.datac(dcifimemload_20),
	.datad(\Selector100~1_combout ),
	.cin(gnd),
	.combout(\Selector96~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector96~1 .lut_mask = 16'hAAAE;
defparam \Selector96~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N12
cycloneive_lcell_comb \Selector97~0 (
// Equation(s):
// \Selector97~0_combout  = (WideOr3 & (dcifimemload_3 & ((!cuifALUSrc_1)))) # (!WideOr3 & (((dcifimemload_9 & cuifALUSrc_1))))

	.dataa(dcifimemload_3),
	.datab(dcifimemload_9),
	.datac(\cu|WideOr3~1_combout ),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector97~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector97~0 .lut_mask = 16'h0CA0;
defparam \Selector97~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N28
cycloneive_lcell_comb \Selector97~1 (
// Equation(s):
// \Selector97~1_combout  = (\Selector97~0_combout ) # ((!dcifimemload_20 & (!\Selector100~1_combout  & Mux601)))

	.dataa(\Selector97~0_combout ),
	.datab(dcifimemload_20),
	.datac(\Selector100~1_combout ),
	.datad(Mux601),
	.cin(gnd),
	.combout(\Selector97~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector97~1 .lut_mask = 16'hABAA;
defparam \Selector97~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N26
cycloneive_lcell_comb \Selector98~0 (
// Equation(s):
// \Selector98~0_combout  = (WideOr3 & (((dcifimemload_2 & !cuifALUSrc_1)))) # (!WideOr3 & (dcifimemload_8 & ((cuifALUSrc_1))))

	.dataa(dcifimemload_8),
	.datab(\cu|WideOr3~1_combout ),
	.datac(dcifimemload_2),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector98~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector98~0 .lut_mask = 16'h22C0;
defparam \Selector98~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N10
cycloneive_lcell_comb \Selector98~1 (
// Equation(s):
// \Selector98~1_combout  = (\Selector98~0_combout ) # ((!\Selector100~1_combout  & (!dcifimemload_20 & Mux611)))

	.dataa(\Selector100~1_combout ),
	.datab(dcifimemload_20),
	.datac(\Selector98~0_combout ),
	.datad(Mux611),
	.cin(gnd),
	.combout(\Selector98~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector98~1 .lut_mask = 16'hF1F0;
defparam \Selector98~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N8
cycloneive_lcell_comb \Selector99~0 (
// Equation(s):
// \Selector99~0_combout  = (WideOr3 & (dcifimemload_1 & ((!cuifALUSrc_1)))) # (!WideOr3 & (((dcifimemload_7 & cuifALUSrc_1))))

	.dataa(dcifimemload_1),
	.datab(dcifimemload_7),
	.datac(\cu|WideOr3~1_combout ),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector99~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector99~0 .lut_mask = 16'h0CA0;
defparam \Selector99~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N10
cycloneive_lcell_comb \Selector99~1 (
// Equation(s):
// \Selector99~1_combout  = (\Selector99~0_combout ) # ((!\Selector100~1_combout  & (!dcifimemload_20 & Mux621)))

	.dataa(\Selector100~1_combout ),
	.datab(dcifimemload_20),
	.datac(\Selector99~0_combout ),
	.datad(Mux621),
	.cin(gnd),
	.combout(\Selector99~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector99~1 .lut_mask = 16'hF1F0;
defparam \Selector99~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N22
cycloneive_lcell_comb \Selector100~2 (
// Equation(s):
// \Selector100~2_combout  = (WideOr3 & (dcifimemload_0 & ((!cuifALUSrc_1)))) # (!WideOr3 & (((dcifimemload_6 & cuifALUSrc_1))))

	.dataa(dcifimemload_0),
	.datab(\cu|WideOr3~1_combout ),
	.datac(dcifimemload_6),
	.datad(\cu|cuif.ALUSrc[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector100~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector100~2 .lut_mask = 16'h3088;
defparam \Selector100~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N28
cycloneive_lcell_comb \Selector100~3 (
// Equation(s):
// \Selector100~3_combout  = (\Selector100~2_combout ) # ((!dcifimemload_20 & (!\Selector100~1_combout  & Mux631)))

	.dataa(dcifimemload_20),
	.datab(\Selector100~1_combout ),
	.datac(\Selector100~2_combout ),
	.datad(Mux631),
	.cin(gnd),
	.combout(\Selector100~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector100~3 .lut_mask = 16'hF1F0;
defparam \Selector100~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N16
cycloneive_lcell_comb \Selector99~2 (
// Equation(s):
// \Selector99~2_combout  = (\Selector99~1_combout ) # ((!\Selector100~1_combout  & (dcifimemload_20 & Mux62)))

	.dataa(\Selector100~1_combout ),
	.datab(dcifimemload_20),
	.datac(Mux62),
	.datad(\Selector99~1_combout ),
	.cin(gnd),
	.combout(\Selector99~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector99~2 .lut_mask = 16'hFF40;
defparam \Selector99~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N30
cycloneive_lcell_comb \Selector100~4 (
// Equation(s):
// \Selector100~4_combout  = (\Selector100~3_combout ) # ((dcifimemload_20 & (Mux63 & !\Selector100~1_combout )))

	.dataa(dcifimemload_20),
	.datab(Mux63),
	.datac(\Selector100~1_combout ),
	.datad(\Selector100~3_combout ),
	.cin(gnd),
	.combout(\Selector100~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector100~4 .lut_mask = 16'hFF08;
defparam \Selector100~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N0
cycloneive_lcell_comb \Selector98~2 (
// Equation(s):
// \Selector98~2_combout  = (\Selector98~1_combout ) # ((!\Selector100~1_combout  & (dcifimemload_20 & Mux61)))

	.dataa(\Selector100~1_combout ),
	.datab(dcifimemload_20),
	.datac(Mux61),
	.datad(\Selector98~1_combout ),
	.cin(gnd),
	.combout(\Selector98~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector98~2 .lut_mask = 16'hFF40;
defparam \Selector98~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N30
cycloneive_lcell_comb \Selector95~3 (
// Equation(s):
// \Selector95~3_combout  = (\Selector95~2_combout ) # ((\Selector95~0_combout  & Mux58))

	.dataa(gnd),
	.datab(\Selector95~0_combout ),
	.datac(Mux58),
	.datad(\Selector95~2_combout ),
	.cin(gnd),
	.combout(\Selector95~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector95~3 .lut_mask = 16'hFFC0;
defparam \Selector95~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N12
cycloneive_lcell_comb \Selector94~1 (
// Equation(s):
// \Selector94~1_combout  = (\Selector94~0_combout ) # ((\Selector95~0_combout  & Mux57))

	.dataa(gnd),
	.datab(\Selector95~0_combout ),
	.datac(\Selector94~0_combout ),
	.datad(Mux57),
	.cin(gnd),
	.combout(\Selector94~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector94~1 .lut_mask = 16'hFCF0;
defparam \Selector94~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N10
cycloneive_lcell_comb \Selector93~1 (
// Equation(s):
// \Selector93~1_combout  = (\Selector93~0_combout ) # ((Mux56 & \Selector95~0_combout ))

	.dataa(Mux56),
	.datab(\Selector95~0_combout ),
	.datac(gnd),
	.datad(\Selector93~0_combout ),
	.cin(gnd),
	.combout(\Selector93~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector93~1 .lut_mask = 16'hFF88;
defparam \Selector93~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N8
cycloneive_lcell_comb \Selector92~1 (
// Equation(s):
// \Selector92~1_combout  = (\Selector92~0_combout ) # ((\Selector95~0_combout  & Mux55))

	.dataa(gnd),
	.datab(\Selector95~0_combout ),
	.datac(Mux55),
	.datad(\Selector92~0_combout ),
	.cin(gnd),
	.combout(\Selector92~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector92~1 .lut_mask = 16'hFFC0;
defparam \Selector92~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N10
cycloneive_lcell_comb \Selector91~1 (
// Equation(s):
// \Selector91~1_combout  = (\Selector91~0_combout ) # ((\Selector95~0_combout  & Mux54))

	.dataa(\Selector95~0_combout ),
	.datab(gnd),
	.datac(Mux54),
	.datad(\Selector91~0_combout ),
	.cin(gnd),
	.combout(\Selector91~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector91~1 .lut_mask = 16'hFFA0;
defparam \Selector91~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N12
cycloneive_lcell_comb \Selector90~1 (
// Equation(s):
// \Selector90~1_combout  = (\Selector90~0_combout ) # ((\Selector95~0_combout  & Mux53))

	.dataa(\Selector95~0_combout ),
	.datab(gnd),
	.datac(\Selector90~0_combout ),
	.datad(Mux53),
	.cin(gnd),
	.combout(\Selector90~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector90~1 .lut_mask = 16'hFAF0;
defparam \Selector90~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N18
cycloneive_lcell_comb \Selector89~1 (
// Equation(s):
// \Selector89~1_combout  = (\Selector89~0_combout ) # ((\Selector95~0_combout  & Mux52))

	.dataa(\Selector95~0_combout ),
	.datab(gnd),
	.datac(\Selector89~0_combout ),
	.datad(Mux52),
	.cin(gnd),
	.combout(\Selector89~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector89~1 .lut_mask = 16'hFAF0;
defparam \Selector89~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N8
cycloneive_lcell_comb \Selector88~1 (
// Equation(s):
// \Selector88~1_combout  = (\Selector88~0_combout ) # ((Mux51 & \Selector95~0_combout ))

	.dataa(Mux51),
	.datab(gnd),
	.datac(\Selector95~0_combout ),
	.datad(\Selector88~0_combout ),
	.cin(gnd),
	.combout(\Selector88~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector88~1 .lut_mask = 16'hFFA0;
defparam \Selector88~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N8
cycloneive_lcell_comb \Selector87~1 (
// Equation(s):
// \Selector87~1_combout  = (\Selector87~0_combout ) # ((Mux50 & \Selector95~0_combout ))

	.dataa(gnd),
	.datab(Mux50),
	.datac(\Selector95~0_combout ),
	.datad(\Selector87~0_combout ),
	.cin(gnd),
	.combout(\Selector87~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector87~1 .lut_mask = 16'hFFC0;
defparam \Selector87~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N24
cycloneive_lcell_comb \Selector86~1 (
// Equation(s):
// \Selector86~1_combout  = (\Selector86~0_combout ) # ((Mux49 & \Selector95~0_combout ))

	.dataa(Mux49),
	.datab(gnd),
	.datac(\Selector95~0_combout ),
	.datad(\Selector86~0_combout ),
	.cin(gnd),
	.combout(\Selector86~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector86~1 .lut_mask = 16'hFFA0;
defparam \Selector86~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N8
cycloneive_lcell_comb \Selector85~1 (
// Equation(s):
// \Selector85~1_combout  = (\Selector85~0_combout ) # ((\Selector95~0_combout  & Mux48))

	.dataa(gnd),
	.datab(\Selector95~0_combout ),
	.datac(\Selector85~0_combout ),
	.datad(Mux48),
	.cin(gnd),
	.combout(\Selector85~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector85~1 .lut_mask = 16'hFCF0;
defparam \Selector85~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N6
cycloneive_lcell_comb \Selector84~2 (
// Equation(s):
// \Selector84~2_combout  = (\Selector84~1_combout ) # ((\Selector95~0_combout  & Mux47))

	.dataa(\Selector95~0_combout ),
	.datab(gnd),
	.datac(Mux47),
	.datad(\Selector84~1_combout ),
	.cin(gnd),
	.combout(\Selector84~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector84~2 .lut_mask = 16'hFFA0;
defparam \Selector84~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N10
cycloneive_lcell_comb \Selector83~1 (
// Equation(s):
// \Selector83~1_combout  = (\Selector83~0_combout ) # ((Mux46 & \Selector95~0_combout ))

	.dataa(Mux46),
	.datab(gnd),
	.datac(\Selector95~0_combout ),
	.datad(\Selector83~0_combout ),
	.cin(gnd),
	.combout(\Selector83~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector83~1 .lut_mask = 16'hFFA0;
defparam \Selector83~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N0
cycloneive_lcell_comb \Selector82~1 (
// Equation(s):
// \Selector82~1_combout  = (\Selector82~0_combout ) # ((\Selector95~0_combout  & Mux45))

	.dataa(\Selector95~0_combout ),
	.datab(gnd),
	.datac(Mux45),
	.datad(\Selector82~0_combout ),
	.cin(gnd),
	.combout(\Selector82~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector82~1 .lut_mask = 16'hFFA0;
defparam \Selector82~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N26
cycloneive_lcell_comb \Selector81~1 (
// Equation(s):
// \Selector81~1_combout  = (\Selector81~0_combout ) # ((Mux44 & \Selector95~0_combout ))

	.dataa(Mux44),
	.datab(gnd),
	.datac(\Selector95~0_combout ),
	.datad(\Selector81~0_combout ),
	.cin(gnd),
	.combout(\Selector81~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector81~1 .lut_mask = 16'hFFA0;
defparam \Selector81~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N4
cycloneive_lcell_comb \Selector80~1 (
// Equation(s):
// \Selector80~1_combout  = (\Selector80~0_combout ) # ((Mux43 & \Selector95~0_combout ))

	.dataa(gnd),
	.datab(Mux43),
	.datac(\Selector95~0_combout ),
	.datad(\Selector80~0_combout ),
	.cin(gnd),
	.combout(\Selector80~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector80~1 .lut_mask = 16'hFFC0;
defparam \Selector80~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N12
cycloneive_lcell_comb \Selector79~1 (
// Equation(s):
// \Selector79~1_combout  = (\Selector79~0_combout ) # ((\Selector95~0_combout  & Mux42))

	.dataa(\Selector95~0_combout ),
	.datab(Mux42),
	.datac(gnd),
	.datad(\Selector79~0_combout ),
	.cin(gnd),
	.combout(\Selector79~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector79~1 .lut_mask = 16'hFF88;
defparam \Selector79~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N20
cycloneive_lcell_comb \Selector78~1 (
// Equation(s):
// \Selector78~1_combout  = (\Selector78~0_combout ) # ((\Selector95~0_combout  & Mux41))

	.dataa(\Selector95~0_combout ),
	.datab(gnd),
	.datac(\Selector78~0_combout ),
	.datad(Mux41),
	.cin(gnd),
	.combout(\Selector78~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector78~1 .lut_mask = 16'hFAF0;
defparam \Selector78~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N26
cycloneive_lcell_comb \Selector77~1 (
// Equation(s):
// \Selector77~1_combout  = (\Selector77~0_combout ) # ((\Selector95~0_combout  & Mux40))

	.dataa(\Selector95~0_combout ),
	.datab(gnd),
	.datac(\Selector77~0_combout ),
	.datad(Mux40),
	.cin(gnd),
	.combout(\Selector77~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector77~1 .lut_mask = 16'hFAF0;
defparam \Selector77~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N0
cycloneive_lcell_comb \Selector76~1 (
// Equation(s):
// \Selector76~1_combout  = (\Selector76~0_combout ) # ((\Selector95~0_combout  & Mux39))

	.dataa(\Selector95~0_combout ),
	.datab(Mux39),
	.datac(\Selector76~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector76~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector76~1 .lut_mask = 16'hF8F8;
defparam \Selector76~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N16
cycloneive_lcell_comb \Selector75~1 (
// Equation(s):
// \Selector75~1_combout  = (\Selector75~0_combout ) # ((Mux38 & \Selector95~0_combout ))

	.dataa(gnd),
	.datab(Mux38),
	.datac(\Selector95~0_combout ),
	.datad(\Selector75~0_combout ),
	.cin(gnd),
	.combout(\Selector75~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector75~1 .lut_mask = 16'hFFC0;
defparam \Selector75~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N18
cycloneive_lcell_comb \Selector74~1 (
// Equation(s):
// \Selector74~1_combout  = (\Selector74~0_combout ) # ((Mux37 & \Selector95~0_combout ))

	.dataa(Mux37),
	.datab(gnd),
	.datac(\Selector95~0_combout ),
	.datad(\Selector74~0_combout ),
	.cin(gnd),
	.combout(\Selector74~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector74~1 .lut_mask = 16'hFFA0;
defparam \Selector74~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N8
cycloneive_lcell_comb \Selector73~1 (
// Equation(s):
// \Selector73~1_combout  = (\Selector73~0_combout ) # ((Mux36 & \Selector95~0_combout ))

	.dataa(Mux36),
	.datab(gnd),
	.datac(\Selector95~0_combout ),
	.datad(\Selector73~0_combout ),
	.cin(gnd),
	.combout(\Selector73~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector73~1 .lut_mask = 16'hFFA0;
defparam \Selector73~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N26
cycloneive_lcell_comb \Selector72~1 (
// Equation(s):
// \Selector72~1_combout  = (\Selector72~0_combout ) # ((Mux35 & \Selector95~0_combout ))

	.dataa(Mux35),
	.datab(gnd),
	.datac(\Selector95~0_combout ),
	.datad(\Selector72~0_combout ),
	.cin(gnd),
	.combout(\Selector72~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector72~1 .lut_mask = 16'hFFA0;
defparam \Selector72~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N6
cycloneive_lcell_comb \Selector71~1 (
// Equation(s):
// \Selector71~1_combout  = (\Selector71~0_combout ) # ((\Selector95~0_combout  & Mux34))

	.dataa(gnd),
	.datab(\Selector71~0_combout ),
	.datac(\Selector95~0_combout ),
	.datad(Mux34),
	.cin(gnd),
	.combout(\Selector71~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector71~1 .lut_mask = 16'hFCCC;
defparam \Selector71~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N30
cycloneive_lcell_comb \Selector70~1 (
// Equation(s):
// \Selector70~1_combout  = (\Selector70~0_combout ) # ((\Selector95~0_combout  & Mux33))

	.dataa(gnd),
	.datab(\Selector95~0_combout ),
	.datac(Mux33),
	.datad(\Selector70~0_combout ),
	.cin(gnd),
	.combout(\Selector70~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector70~1 .lut_mask = 16'hFFC0;
defparam \Selector70~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N18
cycloneive_lcell_comb \Selector69~0 (
// Equation(s):
// \Selector69~0_combout  = (\Selector84~0_combout ) # ((Mux32 & \Selector95~1_combout ))

	.dataa(gnd),
	.datab(Mux32),
	.datac(\Selector95~1_combout ),
	.datad(\Selector84~0_combout ),
	.cin(gnd),
	.combout(\Selector69~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector69~0 .lut_mask = 16'hFFC0;
defparam \Selector69~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N12
cycloneive_lcell_comb \Selector69~1 (
// Equation(s):
// \Selector69~1_combout  = (\Selector69~0_combout ) # ((Mux321 & \Selector95~0_combout ))

	.dataa(gnd),
	.datab(Mux321),
	.datac(\Selector95~0_combout ),
	.datad(\Selector69~0_combout ),
	.cin(gnd),
	.combout(\Selector69~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector69~1 .lut_mask = 16'hFFC0;
defparam \Selector69~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N16
cycloneive_lcell_comb \Selector96~2 (
// Equation(s):
// \Selector96~2_combout  = (\Selector96~1_combout ) # ((\Selector100~0_combout  & Mux59))

	.dataa(gnd),
	.datab(\Selector100~0_combout ),
	.datac(Mux59),
	.datad(\Selector96~1_combout ),
	.cin(gnd),
	.combout(\Selector96~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector96~2 .lut_mask = 16'hFFC0;
defparam \Selector96~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N4
cycloneive_lcell_comb \Selector97~2 (
// Equation(s):
// \Selector97~2_combout  = (\Selector97~1_combout ) # ((Mux60 & \Selector100~0_combout ))

	.dataa(Mux60),
	.datab(gnd),
	.datac(\Selector100~0_combout ),
	.datad(\Selector97~1_combout ),
	.cin(gnd),
	.combout(\Selector97~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector97~2 .lut_mask = 16'hFFA0;
defparam \Selector97~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N14
cycloneive_lcell_comb \Selector68~0 (
// Equation(s):
// \Selector68~0_combout  = (!dcifimemload_30 & ((dcifimemload_29 & (!dcifimemload_31)) # (!dcifimemload_29 & ((Decoder11)))))

	.dataa(dcifimemload_31),
	.datab(dcifimemload_30),
	.datac(\cu|Decoder1~2_combout ),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\Selector68~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector68~0 .lut_mask = 16'h1130;
defparam \Selector68~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N28
cycloneive_lcell_comb \Equal10~0 (
// Equation(s):
// \Equal10~0_combout  = (!dcifimemload_30 & ((dcifimemload_31 & (Decoder11 & !dcifimemload_29)) # (!dcifimemload_31 & ((dcifimemload_29)))))

	.dataa(dcifimemload_31),
	.datab(dcifimemload_30),
	.datac(\cu|Decoder1~2_combout ),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\Equal10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~0 .lut_mask = 16'h1120;
defparam \Equal10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N30
cycloneive_lcell_comb \Selector68~1 (
// Equation(s):
// \Selector68~1_combout  = (dcifimemload_11 & ((dcifimemload_16) # ((!\Equal10~0_combout )))) # (!dcifimemload_11 & (\Selector68~0_combout  & ((dcifimemload_16) # (!\Equal10~0_combout ))))

	.dataa(dcifimemload_11),
	.datab(dcifimemload_16),
	.datac(\Selector68~0_combout ),
	.datad(\Equal10~0_combout ),
	.cin(gnd),
	.combout(\Selector68~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector68~1 .lut_mask = 16'hC8FA;
defparam \Selector68~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N16
cycloneive_lcell_comb \Selector67~0 (
// Equation(s):
// \Selector67~0_combout  = (dcifimemload_12 & ((dcifimemload_17) # ((!\Equal10~0_combout )))) # (!dcifimemload_12 & (\Selector68~0_combout  & ((dcifimemload_17) # (!\Equal10~0_combout ))))

	.dataa(dcifimemload_12),
	.datab(dcifimemload_17),
	.datac(\Selector68~0_combout ),
	.datad(\Equal10~0_combout ),
	.cin(gnd),
	.combout(\Selector67~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector67~0 .lut_mask = 16'hC8FA;
defparam \Selector67~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N20
cycloneive_lcell_comb \Selector64~0 (
// Equation(s):
// \Selector64~0_combout  = (dcifimemload_15 & ((dcifimemload_20) # ((!\Equal10~0_combout )))) # (!dcifimemload_15 & (\Selector68~0_combout  & ((dcifimemload_20) # (!\Equal10~0_combout ))))

	.dataa(dcifimemload_15),
	.datab(dcifimemload_20),
	.datac(\Equal10~0_combout ),
	.datad(\Selector68~0_combout ),
	.cin(gnd),
	.combout(\Selector64~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector64~0 .lut_mask = 16'hCF8A;
defparam \Selector64~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N10
cycloneive_lcell_comb \Selector66~0 (
// Equation(s):
// \Selector66~0_combout  = (dcifimemload_13 & ((dcifimemload_18) # ((!\Equal10~0_combout )))) # (!dcifimemload_13 & (\Selector68~0_combout  & ((dcifimemload_18) # (!\Equal10~0_combout ))))

	.dataa(dcifimemload_13),
	.datab(dcifimemload_18),
	.datac(\Selector68~0_combout ),
	.datad(\Equal10~0_combout ),
	.cin(gnd),
	.combout(\Selector66~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector66~0 .lut_mask = 16'hC8FA;
defparam \Selector66~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N14
cycloneive_lcell_comb \Selector65~0 (
// Equation(s):
// \Selector65~0_combout  = (dcifimemload_14 & ((dcifimemload_19) # ((!\Equal10~0_combout )))) # (!dcifimemload_14 & (\Selector68~0_combout  & ((dcifimemload_19) # (!\Equal10~0_combout ))))

	.dataa(dcifimemload_14),
	.datab(dcifimemload_19),
	.datac(\Equal10~0_combout ),
	.datad(\Selector68~0_combout ),
	.cin(gnd),
	.combout(\Selector65~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector65~0 .lut_mask = 16'hCF8A;
defparam \Selector65~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N0
cycloneive_lcell_comb \Selector1~0 (
// Equation(s):
// \Selector1~0_combout  = (cuifRegSel_11 & (((cuifRegSel_0)))) # (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_301)) # (!cuifRegSel_0 & ((Mux114)))))

	.dataa(ramiframload_30),
	.datab(\cu|cuif.RegSel[1]~5_combout ),
	.datac(\cu|cuif.RegSel[0]~3_combout ),
	.datad(\ALU|Mux1~9_combout ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~0 .lut_mask = 16'hE3E0;
defparam \Selector1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N14
cycloneive_lcell_comb \Selector1~1 (
// Equation(s):
// \Selector1~1_combout  = (cuifRegSel_11 & ((\Selector1~0_combout  & ((dcifimemload_14))) # (!\Selector1~0_combout  & (\Add1~56_combout )))) # (!cuifRegSel_11 & (((\Selector1~0_combout ))))

	.dataa(\Add1~56_combout ),
	.datab(\cu|cuif.RegSel[1]~5_combout ),
	.datac(dcifimemload_14),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~1 .lut_mask = 16'hF388;
defparam \Selector1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N2
cycloneive_lcell_comb \Selector2~0 (
// Equation(s):
// \Selector2~0_combout  = (cuifRegSel_11 & ((\Add1~54_combout ) # ((cuifRegSel_0)))) # (!cuifRegSel_11 & (((!cuifRegSel_0 & Mux210))))

	.dataa(\cu|cuif.RegSel[1]~5_combout ),
	.datab(\Add1~54_combout ),
	.datac(\cu|cuif.RegSel[0]~3_combout ),
	.datad(Mux2),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~0 .lut_mask = 16'hADA8;
defparam \Selector2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N4
cycloneive_lcell_comb \Selector2~1 (
// Equation(s):
// \Selector2~1_combout  = (cuifRegSel_0 & ((\Selector2~0_combout  & (dcifimemload_13)) # (!\Selector2~0_combout  & ((ramiframload_291))))) # (!cuifRegSel_0 & (((\Selector2~0_combout ))))

	.dataa(\cu|cuif.RegSel[0]~3_combout ),
	.datab(dcifimemload_13),
	.datac(ramiframload_29),
	.datad(\Selector2~0_combout ),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~1 .lut_mask = 16'hDDA0;
defparam \Selector2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N10
cycloneive_lcell_comb \Selector3~0 (
// Equation(s):
// \Selector3~0_combout  = (cuifRegSel_0 & ((ramiframload_281) # ((cuifRegSel_11)))) # (!cuifRegSel_0 & (((!cuifRegSel_11 & Mux310))))

	.dataa(\cu|cuif.RegSel[0]~3_combout ),
	.datab(ramiframload_28),
	.datac(\cu|cuif.RegSel[1]~5_combout ),
	.datad(Mux3),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~0 .lut_mask = 16'hADA8;
defparam \Selector3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N28
cycloneive_lcell_comb \Selector3~1 (
// Equation(s):
// \Selector3~1_combout  = (cuifRegSel_11 & ((\Selector3~0_combout  & ((dcifimemload_12))) # (!\Selector3~0_combout  & (\Add1~52_combout )))) # (!cuifRegSel_11 & (((\Selector3~0_combout ))))

	.dataa(\Add1~52_combout ),
	.datab(dcifimemload_12),
	.datac(\cu|cuif.RegSel[1]~5_combout ),
	.datad(\Selector3~0_combout ),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~1 .lut_mask = 16'hCFA0;
defparam \Selector3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N24
cycloneive_lcell_comb \Selector8~0 (
// Equation(s):
// \Selector8~0_combout  = (cuifRegSel_11 & ((\Add1~42_combout ) # ((cuifRegSel_0)))) # (!cuifRegSel_11 & (((!cuifRegSel_0 & Mux81))))

	.dataa(\cu|cuif.RegSel[1]~5_combout ),
	.datab(\Add1~42_combout ),
	.datac(\cu|cuif.RegSel[0]~3_combout ),
	.datad(Mux8),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~0 .lut_mask = 16'hADA8;
defparam \Selector8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N26
cycloneive_lcell_comb \Selector8~1 (
// Equation(s):
// \Selector8~1_combout  = (cuifRegSel_0 & ((\Selector8~0_combout  & ((dcifimemload_7))) # (!\Selector8~0_combout  & (ramiframload_23)))) # (!cuifRegSel_0 & (((\Selector8~0_combout ))))

	.dataa(ramiframload_23),
	.datab(dcifimemload_7),
	.datac(\cu|cuif.RegSel[0]~3_combout ),
	.datad(\Selector8~0_combout ),
	.cin(gnd),
	.combout(\Selector8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~1 .lut_mask = 16'hCFA0;
defparam \Selector8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N28
cycloneive_lcell_comb \Selector9~0 (
// Equation(s):
// \Selector9~0_combout  = (cuifRegSel_0 & ((cuifRegSel_11) # ((ramiframload_22)))) # (!cuifRegSel_0 & (!cuifRegSel_11 & ((Mux93))))

	.dataa(\cu|cuif.RegSel[0]~3_combout ),
	.datab(\cu|cuif.RegSel[1]~5_combout ),
	.datac(ramiframload_22),
	.datad(\ALU|Mux9~9_combout ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~0 .lut_mask = 16'hB9A8;
defparam \Selector9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N26
cycloneive_lcell_comb \Selector9~1 (
// Equation(s):
// \Selector9~1_combout  = (cuifRegSel_11 & ((\Selector9~0_combout  & (dcifimemload_6)) # (!\Selector9~0_combout  & ((\Add1~40_combout ))))) # (!cuifRegSel_11 & (((\Selector9~0_combout ))))

	.dataa(dcifimemload_6),
	.datab(\cu|cuif.RegSel[1]~5_combout ),
	.datac(\Add1~40_combout ),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\Selector9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~1 .lut_mask = 16'hBBC0;
defparam \Selector9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N6
cycloneive_lcell_comb \Selector10~0 (
// Equation(s):
// \Selector10~0_combout  = (cuifRegSel_0 & (((cuifRegSel_11)))) # (!cuifRegSel_0 & ((cuifRegSel_11 & (\Add1~38_combout )) # (!cuifRegSel_11 & ((Mux103)))))

	.dataa(\cu|cuif.RegSel[0]~3_combout ),
	.datab(\Add1~38_combout ),
	.datac(\cu|cuif.RegSel[1]~5_combout ),
	.datad(\ALU|Mux10~7_combout ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~0 .lut_mask = 16'hE5E0;
defparam \Selector10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N8
cycloneive_lcell_comb \Selector10~1 (
// Equation(s):
// \Selector10~1_combout  = (cuifRegSel_0 & ((\Selector10~0_combout  & (dcifimemload_5)) # (!\Selector10~0_combout  & ((ramiframload_211))))) # (!cuifRegSel_0 & (((\Selector10~0_combout ))))

	.dataa(\cu|cuif.RegSel[0]~3_combout ),
	.datab(dcifimemload_5),
	.datac(ramiframload_21),
	.datad(\Selector10~0_combout ),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~1 .lut_mask = 16'hDDA0;
defparam \Selector10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N8
cycloneive_lcell_comb \Selector11~0 (
// Equation(s):
// \Selector11~0_combout  = (cuifRegSel_0 & ((ramiframload_20) # ((cuifRegSel_11)))) # (!cuifRegSel_0 & (((!cuifRegSel_11 & Mux115))))

	.dataa(\cu|cuif.RegSel[0]~3_combout ),
	.datab(ramiframload_20),
	.datac(\cu|cuif.RegSel[1]~5_combout ),
	.datad(\ALU|Mux11~7_combout ),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~0 .lut_mask = 16'hADA8;
defparam \Selector11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N14
cycloneive_lcell_comb \Selector11~1 (
// Equation(s):
// \Selector11~1_combout  = (cuifRegSel_11 & ((\Selector11~0_combout  & (dcifimemload_4)) # (!\Selector11~0_combout  & ((\Add1~36_combout ))))) # (!cuifRegSel_11 & (((\Selector11~0_combout ))))

	.dataa(\cu|cuif.RegSel[1]~5_combout ),
	.datab(dcifimemload_4),
	.datac(\Selector11~0_combout ),
	.datad(\Add1~36_combout ),
	.cin(gnd),
	.combout(\Selector11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~1 .lut_mask = 16'hDAD0;
defparam \Selector11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N2
cycloneive_lcell_comb \Selector12~0 (
// Equation(s):
// \Selector12~0_combout  = (cuifRegSel_11 & ((\Add1~34_combout ) # ((cuifRegSel_0)))) # (!cuifRegSel_11 & (((!cuifRegSel_0 & Mux123))))

	.dataa(\cu|cuif.RegSel[1]~5_combout ),
	.datab(\Add1~34_combout ),
	.datac(\cu|cuif.RegSel[0]~3_combout ),
	.datad(\ALU|Mux12~7_combout ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~0 .lut_mask = 16'hADA8;
defparam \Selector12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N12
cycloneive_lcell_comb \Selector12~1 (
// Equation(s):
// \Selector12~1_combout  = (cuifRegSel_0 & ((\Selector12~0_combout  & (dcifimemload_3)) # (!\Selector12~0_combout  & ((ramiframload_19))))) # (!cuifRegSel_0 & (((\Selector12~0_combout ))))

	.dataa(dcifimemload_3),
	.datab(\cu|cuif.RegSel[0]~3_combout ),
	.datac(ramiframload_19),
	.datad(\Selector12~0_combout ),
	.cin(gnd),
	.combout(\Selector12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~1 .lut_mask = 16'hBBC0;
defparam \Selector12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N28
cycloneive_lcell_comb \Selector13~0 (
// Equation(s):
// \Selector13~0_combout  = (cuifRegSel_0 & ((cuifRegSel_11) # ((ramiframload_18)))) # (!cuifRegSel_0 & (!cuifRegSel_11 & ((Mux133))))

	.dataa(\cu|cuif.RegSel[0]~3_combout ),
	.datab(\cu|cuif.RegSel[1]~5_combout ),
	.datac(ramiframload_18),
	.datad(\ALU|Mux13~7_combout ),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~0 .lut_mask = 16'hB9A8;
defparam \Selector13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N6
cycloneive_lcell_comb \Selector13~1 (
// Equation(s):
// \Selector13~1_combout  = (cuifRegSel_11 & ((\Selector13~0_combout  & (dcifimemload_2)) # (!\Selector13~0_combout  & ((\Add1~32_combout ))))) # (!cuifRegSel_11 & (((\Selector13~0_combout ))))

	.dataa(dcifimemload_2),
	.datab(\cu|cuif.RegSel[1]~5_combout ),
	.datac(\Add1~32_combout ),
	.datad(\Selector13~0_combout ),
	.cin(gnd),
	.combout(\Selector13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~1 .lut_mask = 16'hBBC0;
defparam \Selector13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N28
cycloneive_lcell_comb \Selector14~0 (
// Equation(s):
// \Selector14~0_combout  = (cuifRegSel_0 & (cuifRegSel_11)) # (!cuifRegSel_0 & ((cuifRegSel_11 & (\Add1~30_combout )) # (!cuifRegSel_11 & ((Mux143)))))

	.dataa(\cu|cuif.RegSel[0]~3_combout ),
	.datab(\cu|cuif.RegSel[1]~5_combout ),
	.datac(\Add1~30_combout ),
	.datad(\ALU|Mux14~9_combout ),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~0 .lut_mask = 16'hD9C8;
defparam \Selector14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N0
cycloneive_lcell_comb \Selector14~1 (
// Equation(s):
// \Selector14~1_combout  = (cuifRegSel_0 & ((\Selector14~0_combout  & ((dcifimemload_1))) # (!\Selector14~0_combout  & (ramiframload_171)))) # (!cuifRegSel_0 & (((\Selector14~0_combout ))))

	.dataa(ramiframload_17),
	.datab(dcifimemload_1),
	.datac(\cu|cuif.RegSel[0]~3_combout ),
	.datad(\Selector14~0_combout ),
	.cin(gnd),
	.combout(\Selector14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~1 .lut_mask = 16'hCFA0;
defparam \Selector14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N26
cycloneive_lcell_comb \Selector15~0 (
// Equation(s):
// \Selector15~0_combout  = (cuifRegSel_11 & (((cuifRegSel_0)))) # (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_161)) # (!cuifRegSel_0 & ((Mux153)))))

	.dataa(ramiframload_16),
	.datab(\cu|cuif.RegSel[1]~5_combout ),
	.datac(\cu|cuif.RegSel[0]~3_combout ),
	.datad(\ALU|Mux15~8_combout ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~0 .lut_mask = 16'hE3E0;
defparam \Selector15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N8
cycloneive_lcell_comb \Selector15~1 (
// Equation(s):
// \Selector15~1_combout  = (\Selector15~0_combout  & ((dcifimemload_0) # ((!cuifRegSel_11)))) # (!\Selector15~0_combout  & (((\Add1~28_combout  & cuifRegSel_11))))

	.dataa(\Selector15~0_combout ),
	.datab(dcifimemload_0),
	.datac(\Add1~28_combout ),
	.datad(\cu|cuif.RegSel[1]~5_combout ),
	.cin(gnd),
	.combout(\Selector15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~1 .lut_mask = 16'hD8AA;
defparam \Selector15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N12
cycloneive_lcell_comb \Selector0~0 (
// Equation(s):
// \Selector0~0_combout  = (cuifRegSel_0 & (((cuifRegSel_11)))) # (!cuifRegSel_0 & ((cuifRegSel_11 & (\Add1~58_combout )) # (!cuifRegSel_11 & ((Mux03)))))

	.dataa(\Add1~58_combout ),
	.datab(\cu|cuif.RegSel[0]~3_combout ),
	.datac(\cu|cuif.RegSel[1]~5_combout ),
	.datad(\ALU|Mux0~15_combout ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~0 .lut_mask = 16'hE3E0;
defparam \Selector0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N14
cycloneive_lcell_comb \Selector0~1 (
// Equation(s):
// \Selector0~1_combout  = (cuifRegSel_0 & ((\Selector0~0_combout  & (dcifimemload_15)) # (!\Selector0~0_combout  & ((ramiframload_311))))) # (!cuifRegSel_0 & (((\Selector0~0_combout ))))

	.dataa(dcifimemload_15),
	.datab(ramiframload_31),
	.datac(\cu|cuif.RegSel[0]~3_combout ),
	.datad(\Selector0~0_combout ),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~1 .lut_mask = 16'hAFC0;
defparam \Selector0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N13
dffeas \PC[29] (
	.clk(CLK),
	.d(\PC[29]~1_combout ),
	.asdata(\Add2~54_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(\PC[28]~8_combout ),
	.sload(\cu|Selector6~1_combout ),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_29),
	.prn(vcc));
// synopsys translate_off
defparam \PC[29] .is_wysiwyg = "true";
defparam \PC[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N31
dffeas \PC[28] (
	.clk(CLK),
	.d(\PC[28]~0_combout ),
	.asdata(\Add2~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(\PC[28]~8_combout ),
	.sload(\cu|Selector6~1_combout ),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_28),
	.prn(vcc));
// synopsys translate_off
defparam \PC[28] .is_wysiwyg = "true";
defparam \PC[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N5
dffeas \PC[31] (
	.clk(CLK),
	.d(\PC[31]~3_combout ),
	.asdata(\Add2~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(\PC[28]~8_combout ),
	.sload(\cu|Selector6~1_combout ),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_31),
	.prn(vcc));
// synopsys translate_off
defparam \PC[31] .is_wysiwyg = "true";
defparam \PC[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N23
dffeas \PC[30] (
	.clk(CLK),
	.d(\PC[30]~2_combout ),
	.asdata(\Add2~56_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(\PC[28]~8_combout ),
	.sload(\cu|Selector6~1_combout ),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_30),
	.prn(vcc));
// synopsys translate_off
defparam \PC[30] .is_wysiwyg = "true";
defparam \PC[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N29
dffeas \dpif.halt~_Duplicate_1 (
	.clk(CLK),
	.d(gnd),
	.asdata(\Equal0~1_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dpifhalt),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt~_Duplicate_1 .is_wysiwyg = "true";
defparam \dpif.halt~_Duplicate_1 .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N9
dffeas \PC[1] (
	.clk(CLK),
	.d(\PC[1]~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_1),
	.prn(vcc));
// synopsys translate_off
defparam \PC[1] .is_wysiwyg = "true";
defparam \PC[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N3
dffeas \PC[0] (
	.clk(CLK),
	.d(\PC[0]~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_0),
	.prn(vcc));
// synopsys translate_off
defparam \PC[0] .is_wysiwyg = "true";
defparam \PC[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N9
dffeas \PC[3] (
	.clk(CLK),
	.d(\Selector60~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_3),
	.prn(vcc));
// synopsys translate_off
defparam \PC[3] .is_wysiwyg = "true";
defparam \PC[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N9
dffeas \PC[2] (
	.clk(CLK),
	.d(\Selector61~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_2),
	.prn(vcc));
// synopsys translate_off
defparam \PC[2] .is_wysiwyg = "true";
defparam \PC[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N1
dffeas \PC[5] (
	.clk(CLK),
	.d(\Selector58~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_5),
	.prn(vcc));
// synopsys translate_off
defparam \PC[5] .is_wysiwyg = "true";
defparam \PC[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N29
dffeas \PC[4] (
	.clk(CLK),
	.d(\Selector59~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_4),
	.prn(vcc));
// synopsys translate_off
defparam \PC[4] .is_wysiwyg = "true";
defparam \PC[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N5
dffeas \PC[7] (
	.clk(CLK),
	.d(\Selector56~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_7),
	.prn(vcc));
// synopsys translate_off
defparam \PC[7] .is_wysiwyg = "true";
defparam \PC[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N7
dffeas \PC[6] (
	.clk(CLK),
	.d(\Selector57~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_6),
	.prn(vcc));
// synopsys translate_off
defparam \PC[6] .is_wysiwyg = "true";
defparam \PC[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N27
dffeas \PC[9] (
	.clk(CLK),
	.d(\Selector54~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_9),
	.prn(vcc));
// synopsys translate_off
defparam \PC[9] .is_wysiwyg = "true";
defparam \PC[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N9
dffeas \PC[8] (
	.clk(CLK),
	.d(\Selector55~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_8),
	.prn(vcc));
// synopsys translate_off
defparam \PC[8] .is_wysiwyg = "true";
defparam \PC[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N25
dffeas \PC[11] (
	.clk(CLK),
	.d(\Selector52~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_11),
	.prn(vcc));
// synopsys translate_off
defparam \PC[11] .is_wysiwyg = "true";
defparam \PC[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N27
dffeas \PC[10] (
	.clk(CLK),
	.d(\Selector53~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_10),
	.prn(vcc));
// synopsys translate_off
defparam \PC[10] .is_wysiwyg = "true";
defparam \PC[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N9
dffeas \PC[13] (
	.clk(CLK),
	.d(\Selector50~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_13),
	.prn(vcc));
// synopsys translate_off
defparam \PC[13] .is_wysiwyg = "true";
defparam \PC[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N31
dffeas \PC[12] (
	.clk(CLK),
	.d(\Selector51~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_12),
	.prn(vcc));
// synopsys translate_off
defparam \PC[12] .is_wysiwyg = "true";
defparam \PC[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N13
dffeas \PC[15] (
	.clk(CLK),
	.d(\Selector48~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_15),
	.prn(vcc));
// synopsys translate_off
defparam \PC[15] .is_wysiwyg = "true";
defparam \PC[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N23
dffeas \PC[14] (
	.clk(CLK),
	.d(\Selector49~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_14),
	.prn(vcc));
// synopsys translate_off
defparam \PC[14] .is_wysiwyg = "true";
defparam \PC[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N21
dffeas \PC[17] (
	.clk(CLK),
	.d(\Selector46~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_17),
	.prn(vcc));
// synopsys translate_off
defparam \PC[17] .is_wysiwyg = "true";
defparam \PC[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N31
dffeas \PC[16] (
	.clk(CLK),
	.d(\Selector47~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_16),
	.prn(vcc));
// synopsys translate_off
defparam \PC[16] .is_wysiwyg = "true";
defparam \PC[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N5
dffeas \PC[19] (
	.clk(CLK),
	.d(\Selector44~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_19),
	.prn(vcc));
// synopsys translate_off
defparam \PC[19] .is_wysiwyg = "true";
defparam \PC[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N13
dffeas \PC[18] (
	.clk(CLK),
	.d(\Selector45~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_18),
	.prn(vcc));
// synopsys translate_off
defparam \PC[18] .is_wysiwyg = "true";
defparam \PC[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N5
dffeas \PC[21] (
	.clk(CLK),
	.d(\Selector42~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_21),
	.prn(vcc));
// synopsys translate_off
defparam \PC[21] .is_wysiwyg = "true";
defparam \PC[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N27
dffeas \PC[20] (
	.clk(CLK),
	.d(\Selector43~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_20),
	.prn(vcc));
// synopsys translate_off
defparam \PC[20] .is_wysiwyg = "true";
defparam \PC[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y43_N5
dffeas \PC[23] (
	.clk(CLK),
	.d(\Selector40~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_23),
	.prn(vcc));
// synopsys translate_off
defparam \PC[23] .is_wysiwyg = "true";
defparam \PC[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y43_N31
dffeas \PC[22] (
	.clk(CLK),
	.d(\Selector41~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_22),
	.prn(vcc));
// synopsys translate_off
defparam \PC[22] .is_wysiwyg = "true";
defparam \PC[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N5
dffeas \PC[25] (
	.clk(CLK),
	.d(\Selector38~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_25),
	.prn(vcc));
// synopsys translate_off
defparam \PC[25] .is_wysiwyg = "true";
defparam \PC[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N27
dffeas \PC[24] (
	.clk(CLK),
	.d(\Selector39~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_24),
	.prn(vcc));
// synopsys translate_off
defparam \PC[24] .is_wysiwyg = "true";
defparam \PC[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N27
dffeas \PC[27] (
	.clk(CLK),
	.d(\Selector36~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_27),
	.prn(vcc));
// synopsys translate_off
defparam \PC[27] .is_wysiwyg = "true";
defparam \PC[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N5
dffeas \PC[26] (
	.clk(CLK),
	.d(\Selector37~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_26),
	.prn(vcc));
// synopsys translate_off
defparam \PC[26] .is_wysiwyg = "true";
defparam \PC[26] .power_up = "low";
// synopsys translate_on

// Location: DDIOOUTCELL_X0_Y31_N18
dffeas \dpif.halt (
	.clk(CLK),
	.d(\Equal0~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dpif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dpifhalt1),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt .is_wysiwyg = "true";
defparam \dpif.halt .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N2
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = PC_2 $ (VCC)
// \Add1~1  = CARRY(PC_2)

	.dataa(PC_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h55AA;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N4
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (PC_3 & (!\Add1~1 )) # (!PC_3 & ((\Add1~1 ) # (GND)))
// \Add1~3  = CARRY((!\Add1~1 ) # (!PC_3))

	.dataa(PC_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h5A5F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N6
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = (PC_4 & (\Add1~3  $ (GND))) # (!PC_4 & (!\Add1~3  & VCC))
// \Add1~5  = CARRY((PC_4 & !\Add1~3 ))

	.dataa(PC_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hA50A;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N8
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (PC_5 & (!\Add1~5 )) # (!PC_5 & ((\Add1~5 ) # (GND)))
// \Add1~7  = CARRY((!\Add1~5 ) # (!PC_5))

	.dataa(gnd),
	.datab(PC_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h3C3F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N10
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = (PC_6 & (\Add1~7  $ (GND))) # (!PC_6 & (!\Add1~7  & VCC))
// \Add1~9  = CARRY((PC_6 & !\Add1~7 ))

	.dataa(gnd),
	.datab(PC_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N12
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (PC_7 & (!\Add1~9 )) # (!PC_7 & ((\Add1~9 ) # (GND)))
// \Add1~11  = CARRY((!\Add1~9 ) # (!PC_7))

	.dataa(gnd),
	.datab(PC_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h3C3F;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N14
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = (PC_8 & (\Add1~11  $ (GND))) # (!PC_8 & (!\Add1~11  & VCC))
// \Add1~13  = CARRY((PC_8 & !\Add1~11 ))

	.dataa(PC_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'hA50A;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N16
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (PC_9 & (!\Add1~13 )) # (!PC_9 & ((\Add1~13 ) # (GND)))
// \Add1~15  = CARRY((!\Add1~13 ) # (!PC_9))

	.dataa(gnd),
	.datab(PC_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h3C3F;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N18
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = (PC_10 & (\Add1~15  $ (GND))) # (!PC_10 & (!\Add1~15  & VCC))
// \Add1~17  = CARRY((PC_10 & !\Add1~15 ))

	.dataa(PC_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'hA50A;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N22
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = (PC_12 & (\Add1~19  $ (GND))) # (!PC_12 & (!\Add1~19  & VCC))
// \Add1~21  = CARRY((PC_12 & !\Add1~19 ))

	.dataa(PC_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'hA50A;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N24
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (PC_13 & (!\Add1~21 )) # (!PC_13 & ((\Add1~21 ) # (GND)))
// \Add1~23  = CARRY((!\Add1~21 ) # (!PC_13))

	.dataa(gnd),
	.datab(PC_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h3C3F;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N26
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = (PC_14 & (\Add1~23  $ (GND))) # (!PC_14 & (!\Add1~23  & VCC))
// \Add1~25  = CARRY((PC_14 & !\Add1~23 ))

	.dataa(PC_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'hA50A;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N28
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (PC_15 & (!\Add1~25 )) # (!PC_15 & ((\Add1~25 ) # (GND)))
// \Add1~27  = CARRY((!\Add1~25 ) # (!PC_15))

	.dataa(gnd),
	.datab(PC_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h3C3F;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N30
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = (PC_16 & (\Add1~27  $ (GND))) # (!PC_16 & (!\Add1~27  & VCC))
// \Add1~29  = CARRY((PC_16 & !\Add1~27 ))

	.dataa(PC_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'hA50A;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N0
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (PC_17 & (!\Add1~29 )) # (!PC_17 & ((\Add1~29 ) # (GND)))
// \Add1~31  = CARRY((!\Add1~29 ) # (!PC_17))

	.dataa(PC_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h5A5F;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N2
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = (PC_18 & (\Add1~31  $ (GND))) # (!PC_18 & (!\Add1~31  & VCC))
// \Add1~33  = CARRY((PC_18 & !\Add1~31 ))

	.dataa(PC_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'hA50A;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N4
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (PC_19 & (!\Add1~33 )) # (!PC_19 & ((\Add1~33 ) # (GND)))
// \Add1~35  = CARRY((!\Add1~33 ) # (!PC_19))

	.dataa(PC_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h5A5F;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N6
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = (PC_20 & (\Add1~35  $ (GND))) # (!PC_20 & (!\Add1~35  & VCC))
// \Add1~37  = CARRY((PC_20 & !\Add1~35 ))

	.dataa(gnd),
	.datab(PC_20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'hC30C;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N8
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (PC_21 & (!\Add1~37 )) # (!PC_21 & ((\Add1~37 ) # (GND)))
// \Add1~39  = CARRY((!\Add1~37 ) # (!PC_21))

	.dataa(PC_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h5A5F;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N10
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = (PC_22 & (\Add1~39  $ (GND))) # (!PC_22 & (!\Add1~39  & VCC))
// \Add1~41  = CARRY((PC_22 & !\Add1~39 ))

	.dataa(gnd),
	.datab(PC_22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'hC30C;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N12
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (PC_23 & (!\Add1~41 )) # (!PC_23 & ((\Add1~41 ) # (GND)))
// \Add1~43  = CARRY((!\Add1~41 ) # (!PC_23))

	.dataa(PC_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h5A5F;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N16
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (PC_25 & (!\Add1~45 )) # (!PC_25 & ((\Add1~45 ) # (GND)))
// \Add1~47  = CARRY((!\Add1~45 ) # (!PC_25))

	.dataa(PC_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h5A5F;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N22
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = (PC_28 & (\Add1~51  $ (GND))) # (!PC_28 & (!\Add1~51  & VCC))
// \Add1~53  = CARRY((PC_28 & !\Add1~51 ))

	.dataa(gnd),
	.datab(PC_28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'hC30C;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N24
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (PC_29 & (!\Add1~53 )) # (!PC_29 & ((\Add1~53 ) # (GND)))
// \Add1~55  = CARRY((!\Add1~53 ) # (!PC_29))

	.dataa(gnd),
	.datab(PC_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h3C3F;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N12
cycloneive_lcell_comb \PC[29]~1 (
// Equation(s):
// \PC[29]~1_combout  = (Selector5 & (Mux2)) # (!Selector5 & ((\Add1~54_combout )))

	.dataa(\rf|Mux2~20_combout ),
	.datab(\cu|Selector5~2_combout ),
	.datac(gnd),
	.datad(\Add1~54_combout ),
	.cin(gnd),
	.combout(\PC[29]~1_combout ),
	.cout());
// synopsys translate_off
defparam \PC[29]~1 .lut_mask = 16'hBB88;
defparam \PC[29]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N2
cycloneive_lcell_comb \Add2~0 (
// Equation(s):
// \Add2~0_combout  = (dcifimemload_0 & (\Add1~0_combout  $ (VCC))) # (!dcifimemload_0 & (\Add1~0_combout  & VCC))
// \Add2~1  = CARRY((dcifimemload_0 & \Add1~0_combout ))

	.dataa(dcifimemload_0),
	.datab(\Add1~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
// synopsys translate_off
defparam \Add2~0 .lut_mask = 16'h6688;
defparam \Add2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N4
cycloneive_lcell_comb \Add2~2 (
// Equation(s):
// \Add2~2_combout  = (\Add1~2_combout  & ((dcifimemload_1 & (\Add2~1  & VCC)) # (!dcifimemload_1 & (!\Add2~1 )))) # (!\Add1~2_combout  & ((dcifimemload_1 & (!\Add2~1 )) # (!dcifimemload_1 & ((\Add2~1 ) # (GND)))))
// \Add2~3  = CARRY((\Add1~2_combout  & (!dcifimemload_1 & !\Add2~1 )) # (!\Add1~2_combout  & ((!\Add2~1 ) # (!dcifimemload_1))))

	.dataa(\Add1~2_combout ),
	.datab(dcifimemload_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
// synopsys translate_off
defparam \Add2~2 .lut_mask = 16'h9617;
defparam \Add2~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N6
cycloneive_lcell_comb \Add2~4 (
// Equation(s):
// \Add2~4_combout  = ((dcifimemload_2 $ (\Add1~4_combout  $ (!\Add2~3 )))) # (GND)
// \Add2~5  = CARRY((dcifimemload_2 & ((\Add1~4_combout ) # (!\Add2~3 ))) # (!dcifimemload_2 & (\Add1~4_combout  & !\Add2~3 )))

	.dataa(dcifimemload_2),
	.datab(\Add1~4_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
// synopsys translate_off
defparam \Add2~4 .lut_mask = 16'h698E;
defparam \Add2~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N8
cycloneive_lcell_comb \Add2~6 (
// Equation(s):
// \Add2~6_combout  = (dcifimemload_3 & ((\Add1~6_combout  & (\Add2~5  & VCC)) # (!\Add1~6_combout  & (!\Add2~5 )))) # (!dcifimemload_3 & ((\Add1~6_combout  & (!\Add2~5 )) # (!\Add1~6_combout  & ((\Add2~5 ) # (GND)))))
// \Add2~7  = CARRY((dcifimemload_3 & (!\Add1~6_combout  & !\Add2~5 )) # (!dcifimemload_3 & ((!\Add2~5 ) # (!\Add1~6_combout ))))

	.dataa(dcifimemload_3),
	.datab(\Add1~6_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
// synopsys translate_off
defparam \Add2~6 .lut_mask = 16'h9617;
defparam \Add2~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N12
cycloneive_lcell_comb \Add2~10 (
// Equation(s):
// \Add2~10_combout  = (dcifimemload_5 & ((\Add1~10_combout  & (\Add2~9  & VCC)) # (!\Add1~10_combout  & (!\Add2~9 )))) # (!dcifimemload_5 & ((\Add1~10_combout  & (!\Add2~9 )) # (!\Add1~10_combout  & ((\Add2~9 ) # (GND)))))
// \Add2~11  = CARRY((dcifimemload_5 & (!\Add1~10_combout  & !\Add2~9 )) # (!dcifimemload_5 & ((!\Add2~9 ) # (!\Add1~10_combout ))))

	.dataa(dcifimemload_5),
	.datab(\Add1~10_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~9 ),
	.combout(\Add2~10_combout ),
	.cout(\Add2~11 ));
// synopsys translate_off
defparam \Add2~10 .lut_mask = 16'h9617;
defparam \Add2~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N14
cycloneive_lcell_comb \Add2~12 (
// Equation(s):
// \Add2~12_combout  = ((dcifimemload_6 $ (\Add1~12_combout  $ (!\Add2~11 )))) # (GND)
// \Add2~13  = CARRY((dcifimemload_6 & ((\Add1~12_combout ) # (!\Add2~11 ))) # (!dcifimemload_6 & (\Add1~12_combout  & !\Add2~11 )))

	.dataa(dcifimemload_6),
	.datab(\Add1~12_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~11 ),
	.combout(\Add2~12_combout ),
	.cout(\Add2~13 ));
// synopsys translate_off
defparam \Add2~12 .lut_mask = 16'h698E;
defparam \Add2~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N16
cycloneive_lcell_comb \Add2~14 (
// Equation(s):
// \Add2~14_combout  = (dcifimemload_7 & ((\Add1~14_combout  & (\Add2~13  & VCC)) # (!\Add1~14_combout  & (!\Add2~13 )))) # (!dcifimemload_7 & ((\Add1~14_combout  & (!\Add2~13 )) # (!\Add1~14_combout  & ((\Add2~13 ) # (GND)))))
// \Add2~15  = CARRY((dcifimemload_7 & (!\Add1~14_combout  & !\Add2~13 )) # (!dcifimemload_7 & ((!\Add2~13 ) # (!\Add1~14_combout ))))

	.dataa(dcifimemload_7),
	.datab(\Add1~14_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~13 ),
	.combout(\Add2~14_combout ),
	.cout(\Add2~15 ));
// synopsys translate_off
defparam \Add2~14 .lut_mask = 16'h9617;
defparam \Add2~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N20
cycloneive_lcell_comb \Add2~18 (
// Equation(s):
// \Add2~18_combout  = (\Add1~18_combout  & ((dcifimemload_9 & (\Add2~17  & VCC)) # (!dcifimemload_9 & (!\Add2~17 )))) # (!\Add1~18_combout  & ((dcifimemload_9 & (!\Add2~17 )) # (!dcifimemload_9 & ((\Add2~17 ) # (GND)))))
// \Add2~19  = CARRY((\Add1~18_combout  & (!dcifimemload_9 & !\Add2~17 )) # (!\Add1~18_combout  & ((!\Add2~17 ) # (!dcifimemload_9))))

	.dataa(\Add1~18_combout ),
	.datab(dcifimemload_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~17 ),
	.combout(\Add2~18_combout ),
	.cout(\Add2~19 ));
// synopsys translate_off
defparam \Add2~18 .lut_mask = 16'h9617;
defparam \Add2~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N22
cycloneive_lcell_comb \Add2~20 (
// Equation(s):
// \Add2~20_combout  = ((dcifimemload_10 $ (\Add1~20_combout  $ (!\Add2~19 )))) # (GND)
// \Add2~21  = CARRY((dcifimemload_10 & ((\Add1~20_combout ) # (!\Add2~19 ))) # (!dcifimemload_10 & (\Add1~20_combout  & !\Add2~19 )))

	.dataa(dcifimemload_10),
	.datab(\Add1~20_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~19 ),
	.combout(\Add2~20_combout ),
	.cout(\Add2~21 ));
// synopsys translate_off
defparam \Add2~20 .lut_mask = 16'h698E;
defparam \Add2~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N24
cycloneive_lcell_comb \Add2~22 (
// Equation(s):
// \Add2~22_combout  = (dcifimemload_11 & ((\Add1~22_combout  & (\Add2~21  & VCC)) # (!\Add1~22_combout  & (!\Add2~21 )))) # (!dcifimemload_11 & ((\Add1~22_combout  & (!\Add2~21 )) # (!\Add1~22_combout  & ((\Add2~21 ) # (GND)))))
// \Add2~23  = CARRY((dcifimemload_11 & (!\Add1~22_combout  & !\Add2~21 )) # (!dcifimemload_11 & ((!\Add2~21 ) # (!\Add1~22_combout ))))

	.dataa(dcifimemload_11),
	.datab(\Add1~22_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~21 ),
	.combout(\Add2~22_combout ),
	.cout(\Add2~23 ));
// synopsys translate_off
defparam \Add2~22 .lut_mask = 16'h9617;
defparam \Add2~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N28
cycloneive_lcell_comb \Add2~26 (
// Equation(s):
// \Add2~26_combout  = (dcifimemload_13 & ((\Add1~26_combout  & (\Add2~25  & VCC)) # (!\Add1~26_combout  & (!\Add2~25 )))) # (!dcifimemload_13 & ((\Add1~26_combout  & (!\Add2~25 )) # (!\Add1~26_combout  & ((\Add2~25 ) # (GND)))))
// \Add2~27  = CARRY((dcifimemload_13 & (!\Add1~26_combout  & !\Add2~25 )) # (!dcifimemload_13 & ((!\Add2~25 ) # (!\Add1~26_combout ))))

	.dataa(dcifimemload_13),
	.datab(\Add1~26_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~25 ),
	.combout(\Add2~26_combout ),
	.cout(\Add2~27 ));
// synopsys translate_off
defparam \Add2~26 .lut_mask = 16'h9617;
defparam \Add2~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N30
cycloneive_lcell_comb \Add2~28 (
// Equation(s):
// \Add2~28_combout  = ((\Add1~28_combout  $ (dcifimemload_14 $ (!\Add2~27 )))) # (GND)
// \Add2~29  = CARRY((\Add1~28_combout  & ((dcifimemload_14) # (!\Add2~27 ))) # (!\Add1~28_combout  & (dcifimemload_14 & !\Add2~27 )))

	.dataa(\Add1~28_combout ),
	.datab(dcifimemload_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~27 ),
	.combout(\Add2~28_combout ),
	.cout(\Add2~29 ));
// synopsys translate_off
defparam \Add2~28 .lut_mask = 16'h698E;
defparam \Add2~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N0
cycloneive_lcell_comb \Add2~30 (
// Equation(s):
// \Add2~30_combout  = (dcifimemload_15 & ((\Add1~30_combout  & (\Add2~29  & VCC)) # (!\Add1~30_combout  & (!\Add2~29 )))) # (!dcifimemload_15 & ((\Add1~30_combout  & (!\Add2~29 )) # (!\Add1~30_combout  & ((\Add2~29 ) # (GND)))))
// \Add2~31  = CARRY((dcifimemload_15 & (!\Add1~30_combout  & !\Add2~29 )) # (!dcifimemload_15 & ((!\Add2~29 ) # (!\Add1~30_combout ))))

	.dataa(dcifimemload_15),
	.datab(\Add1~30_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~29 ),
	.combout(\Add2~30_combout ),
	.cout(\Add2~31 ));
// synopsys translate_off
defparam \Add2~30 .lut_mask = 16'h9617;
defparam \Add2~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N4
cycloneive_lcell_comb \Add2~34 (
// Equation(s):
// \Add2~34_combout  = (dcifimemload_15 & ((\Add1~34_combout  & (\Add2~33  & VCC)) # (!\Add1~34_combout  & (!\Add2~33 )))) # (!dcifimemload_15 & ((\Add1~34_combout  & (!\Add2~33 )) # (!\Add1~34_combout  & ((\Add2~33 ) # (GND)))))
// \Add2~35  = CARRY((dcifimemload_15 & (!\Add1~34_combout  & !\Add2~33 )) # (!dcifimemload_15 & ((!\Add2~33 ) # (!\Add1~34_combout ))))

	.dataa(dcifimemload_15),
	.datab(\Add1~34_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~33 ),
	.combout(\Add2~34_combout ),
	.cout(\Add2~35 ));
// synopsys translate_off
defparam \Add2~34 .lut_mask = 16'h9617;
defparam \Add2~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N6
cycloneive_lcell_comb \Add2~36 (
// Equation(s):
// \Add2~36_combout  = ((dcifimemload_15 $ (\Add1~36_combout  $ (!\Add2~35 )))) # (GND)
// \Add2~37  = CARRY((dcifimemload_15 & ((\Add1~36_combout ) # (!\Add2~35 ))) # (!dcifimemload_15 & (\Add1~36_combout  & !\Add2~35 )))

	.dataa(dcifimemload_15),
	.datab(\Add1~36_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~35 ),
	.combout(\Add2~36_combout ),
	.cout(\Add2~37 ));
// synopsys translate_off
defparam \Add2~36 .lut_mask = 16'h698E;
defparam \Add2~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N8
cycloneive_lcell_comb \Add2~38 (
// Equation(s):
// \Add2~38_combout  = (dcifimemload_15 & ((\Add1~38_combout  & (\Add2~37  & VCC)) # (!\Add1~38_combout  & (!\Add2~37 )))) # (!dcifimemload_15 & ((\Add1~38_combout  & (!\Add2~37 )) # (!\Add1~38_combout  & ((\Add2~37 ) # (GND)))))
// \Add2~39  = CARRY((dcifimemload_15 & (!\Add1~38_combout  & !\Add2~37 )) # (!dcifimemload_15 & ((!\Add2~37 ) # (!\Add1~38_combout ))))

	.dataa(dcifimemload_15),
	.datab(\Add1~38_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~37 ),
	.combout(\Add2~38_combout ),
	.cout(\Add2~39 ));
// synopsys translate_off
defparam \Add2~38 .lut_mask = 16'h9617;
defparam \Add2~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N12
cycloneive_lcell_comb \Add2~42 (
// Equation(s):
// \Add2~42_combout  = (dcifimemload_15 & ((\Add1~42_combout  & (\Add2~41  & VCC)) # (!\Add1~42_combout  & (!\Add2~41 )))) # (!dcifimemload_15 & ((\Add1~42_combout  & (!\Add2~41 )) # (!\Add1~42_combout  & ((\Add2~41 ) # (GND)))))
// \Add2~43  = CARRY((dcifimemload_15 & (!\Add1~42_combout  & !\Add2~41 )) # (!dcifimemload_15 & ((!\Add2~41 ) # (!\Add1~42_combout ))))

	.dataa(dcifimemload_15),
	.datab(\Add1~42_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~41 ),
	.combout(\Add2~42_combout ),
	.cout(\Add2~43 ));
// synopsys translate_off
defparam \Add2~42 .lut_mask = 16'h9617;
defparam \Add2~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N14
cycloneive_lcell_comb \Add2~44 (
// Equation(s):
// \Add2~44_combout  = ((\Add1~44_combout  $ (dcifimemload_15 $ (!\Add2~43 )))) # (GND)
// \Add2~45  = CARRY((\Add1~44_combout  & ((dcifimemload_15) # (!\Add2~43 ))) # (!\Add1~44_combout  & (dcifimemload_15 & !\Add2~43 )))

	.dataa(\Add1~44_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~43 ),
	.combout(\Add2~44_combout ),
	.cout(\Add2~45 ));
// synopsys translate_off
defparam \Add2~44 .lut_mask = 16'h698E;
defparam \Add2~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N16
cycloneive_lcell_comb \Add2~46 (
// Equation(s):
// \Add2~46_combout  = (\Add1~46_combout  & ((dcifimemload_15 & (\Add2~45  & VCC)) # (!dcifimemload_15 & (!\Add2~45 )))) # (!\Add1~46_combout  & ((dcifimemload_15 & (!\Add2~45 )) # (!dcifimemload_15 & ((\Add2~45 ) # (GND)))))
// \Add2~47  = CARRY((\Add1~46_combout  & (!dcifimemload_15 & !\Add2~45 )) # (!\Add1~46_combout  & ((!\Add2~45 ) # (!dcifimemload_15))))

	.dataa(\Add1~46_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~45 ),
	.combout(\Add2~46_combout ),
	.cout(\Add2~47 ));
// synopsys translate_off
defparam \Add2~46 .lut_mask = 16'h9617;
defparam \Add2~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N18
cycloneive_lcell_comb \Add2~48 (
// Equation(s):
// \Add2~48_combout  = ((\Add1~48_combout  $ (dcifimemload_15 $ (!\Add2~47 )))) # (GND)
// \Add2~49  = CARRY((\Add1~48_combout  & ((dcifimemload_15) # (!\Add2~47 ))) # (!\Add1~48_combout  & (dcifimemload_15 & !\Add2~47 )))

	.dataa(\Add1~48_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~47 ),
	.combout(\Add2~48_combout ),
	.cout(\Add2~49 ));
// synopsys translate_off
defparam \Add2~48 .lut_mask = 16'h698E;
defparam \Add2~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N20
cycloneive_lcell_comb \Add2~50 (
// Equation(s):
// \Add2~50_combout  = (\Add1~50_combout  & ((dcifimemload_15 & (\Add2~49  & VCC)) # (!dcifimemload_15 & (!\Add2~49 )))) # (!\Add1~50_combout  & ((dcifimemload_15 & (!\Add2~49 )) # (!dcifimemload_15 & ((\Add2~49 ) # (GND)))))
// \Add2~51  = CARRY((\Add1~50_combout  & (!dcifimemload_15 & !\Add2~49 )) # (!\Add1~50_combout  & ((!\Add2~49 ) # (!dcifimemload_15))))

	.dataa(\Add1~50_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~49 ),
	.combout(\Add2~50_combout ),
	.cout(\Add2~51 ));
// synopsys translate_off
defparam \Add2~50 .lut_mask = 16'h9617;
defparam \Add2~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N22
cycloneive_lcell_comb \Add2~52 (
// Equation(s):
// \Add2~52_combout  = ((\Add1~52_combout  $ (dcifimemload_15 $ (!\Add2~51 )))) # (GND)
// \Add2~53  = CARRY((\Add1~52_combout  & ((dcifimemload_15) # (!\Add2~51 ))) # (!\Add1~52_combout  & (dcifimemload_15 & !\Add2~51 )))

	.dataa(\Add1~52_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~51 ),
	.combout(\Add2~52_combout ),
	.cout(\Add2~53 ));
// synopsys translate_off
defparam \Add2~52 .lut_mask = 16'h698E;
defparam \Add2~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N24
cycloneive_lcell_comb \Add2~54 (
// Equation(s):
// \Add2~54_combout  = (\Add1~54_combout  & ((dcifimemload_15 & (\Add2~53  & VCC)) # (!dcifimemload_15 & (!\Add2~53 )))) # (!\Add1~54_combout  & ((dcifimemload_15 & (!\Add2~53 )) # (!dcifimemload_15 & ((\Add2~53 ) # (GND)))))
// \Add2~55  = CARRY((\Add1~54_combout  & (!dcifimemload_15 & !\Add2~53 )) # (!\Add1~54_combout  & ((!\Add2~53 ) # (!dcifimemload_15))))

	.dataa(\Add1~54_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~53 ),
	.combout(\Add2~54_combout ),
	.cout(\Add2~55 ));
// synopsys translate_off
defparam \Add2~54 .lut_mask = 16'h9617;
defparam \Add2~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N16
cycloneive_lcell_comb \PC[28]~8 (
// Equation(s):
// \PC[28]~8_combout  = (Selector5 & Selector6)

	.dataa(\cu|Selector5~2_combout ),
	.datab(gnd),
	.datac(\cu|Selector6~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\PC[28]~8_combout ),
	.cout());
// synopsys translate_off
defparam \PC[28]~8 .lut_mask = 16'hA0A0;
defparam \PC[28]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N30
cycloneive_lcell_comb \PC[28]~0 (
// Equation(s):
// \PC[28]~0_combout  = (Selector5 & (Mux3)) # (!Selector5 & ((\Add1~52_combout )))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\rf|Mux3~20_combout ),
	.datac(gnd),
	.datad(\Add1~52_combout ),
	.cin(gnd),
	.combout(\PC[28]~0_combout ),
	.cout());
// synopsys translate_off
defparam \PC[28]~0 .lut_mask = 16'hDD88;
defparam \PC[28]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N26
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = (PC_30 & (\Add1~55  $ (GND))) # (!PC_30 & (!\Add1~55  & VCC))
// \Add1~57  = CARRY((PC_30 & !\Add1~55 ))

	.dataa(PC_30),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'hA50A;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N28
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = \Add1~57  $ (PC_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(PC_31),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'h0FF0;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N4
cycloneive_lcell_comb \PC[31]~3 (
// Equation(s):
// \PC[31]~3_combout  = (Selector5 & (Mux0)) # (!Selector5 & ((\Add1~58_combout )))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\rf|Mux0~20_combout ),
	.datac(gnd),
	.datad(\Add1~58_combout ),
	.cin(gnd),
	.combout(\PC[31]~3_combout ),
	.cout());
// synopsys translate_off
defparam \PC[31]~3 .lut_mask = 16'hDD88;
defparam \PC[31]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N26
cycloneive_lcell_comb \Add2~56 (
// Equation(s):
// \Add2~56_combout  = ((\Add1~56_combout  $ (dcifimemload_15 $ (!\Add2~55 )))) # (GND)
// \Add2~57  = CARRY((\Add1~56_combout  & ((dcifimemload_15) # (!\Add2~55 ))) # (!\Add1~56_combout  & (dcifimemload_15 & !\Add2~55 )))

	.dataa(\Add1~56_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~55 ),
	.combout(\Add2~56_combout ),
	.cout(\Add2~57 ));
// synopsys translate_off
defparam \Add2~56 .lut_mask = 16'h698E;
defparam \Add2~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N28
cycloneive_lcell_comb \Add2~58 (
// Equation(s):
// \Add2~58_combout  = dcifimemload_15 $ (\Add1~58_combout  $ (\Add2~57 ))

	.dataa(dcifimemload_15),
	.datab(\Add1~58_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add2~57 ),
	.combout(\Add2~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add2~58 .lut_mask = 16'h9696;
defparam \Add2~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N22
cycloneive_lcell_comb \PC[30]~2 (
// Equation(s):
// \PC[30]~2_combout  = (Selector5 & (Mux1)) # (!Selector5 & ((\Add1~56_combout )))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\rf|Mux1~20_combout ),
	.datac(gnd),
	.datad(\Add1~56_combout ),
	.cin(gnd),
	.combout(\PC[30]~2_combout ),
	.cout());
// synopsys translate_off
defparam \PC[30]~2 .lut_mask = 16'hDD88;
defparam \PC[30]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N16
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (dcifimemload_28 & (dcifimemload_29 & (dcifimemload_30 & dcifimemload_31)))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_29),
	.datac(dcifimemload_30),
	.datad(dcifimemload_31),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h8000;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N12
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// \Equal0~1_combout  = (dcifimemload_27 & (dcifimemload_26 & \Equal0~0_combout ))

	.dataa(dcifimemload_27),
	.datab(gnd),
	.datac(dcifimemload_26),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'hA000;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N0
cycloneive_lcell_comb \PC[0]~9 (
// Equation(s):
// \PC[0]~9_combout  = (Selector5 & (!ccifiwait_01 & !dpifhalt))

	.dataa(\cu|Selector5~2_combout ),
	.datab(ccifiwait_01),
	.datac(gnd),
	.datad(dpifhalt),
	.cin(gnd),
	.combout(\PC[0]~9_combout ),
	.cout());
// synopsys translate_off
defparam \PC[0]~9 .lut_mask = 16'h0022;
defparam \PC[0]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N8
cycloneive_lcell_comb \PC[1]~6 (
// Equation(s):
// \PC[1]~6_combout  = (\PC[0]~9_combout  & (Mux30 & ((!Selector6)))) # (!\PC[0]~9_combout  & (((PC_1))))

	.dataa(\rf|Mux30~20_combout ),
	.datab(\PC[0]~9_combout ),
	.datac(PC_1),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\PC[1]~6_combout ),
	.cout());
// synopsys translate_off
defparam \PC[1]~6 .lut_mask = 16'h30B8;
defparam \PC[1]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N2
cycloneive_lcell_comb \PC[0]~7 (
// Equation(s):
// \PC[0]~7_combout  = (\PC[0]~9_combout  & (Mux31 & ((!Selector6)))) # (!\PC[0]~9_combout  & (((PC_0))))

	.dataa(\PC[0]~9_combout ),
	.datab(\rf|Mux31~20_combout ),
	.datac(PC_0),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\PC[0]~7_combout ),
	.cout());
// synopsys translate_off
defparam \PC[0]~7 .lut_mask = 16'h50D8;
defparam \PC[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N30
cycloneive_lcell_comb \Selector60~0 (
// Equation(s):
// \Selector60~0_combout  = (Selector6 & (((Selector5)))) # (!Selector6 & ((Selector5 & (Mux28)) # (!Selector5 & ((\Add1~2_combout )))))

	.dataa(\rf|Mux28~20_combout ),
	.datab(\Add1~2_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\cu|Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector60~0 .lut_mask = 16'hFA0C;
defparam \Selector60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N8
cycloneive_lcell_comb \Selector60~1 (
// Equation(s):
// \Selector60~1_combout  = (Selector6 & ((\Selector60~0_combout  & (dcifimemload_1)) # (!\Selector60~0_combout  & ((\Add2~2_combout ))))) # (!Selector6 & (((\Selector60~0_combout ))))

	.dataa(\cu|Selector6~1_combout ),
	.datab(dcifimemload_1),
	.datac(\Selector60~0_combout ),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Selector60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector60~1 .lut_mask = 16'hDAD0;
defparam \Selector60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N12
cycloneive_lcell_comb \Selector61~0 (
// Equation(s):
// \Selector61~0_combout  = (Selector6 & ((Selector5) # ((\Add2~0_combout )))) # (!Selector6 & (!Selector5 & (\Add1~0_combout )))

	.dataa(\cu|Selector6~1_combout ),
	.datab(\cu|Selector5~2_combout ),
	.datac(\Add1~0_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Selector61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector61~0 .lut_mask = 16'hBA98;
defparam \Selector61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N8
cycloneive_lcell_comb \Selector61~1 (
// Equation(s):
// \Selector61~1_combout  = (Selector5 & ((\Selector61~0_combout  & ((dcifimemload_0))) # (!\Selector61~0_combout  & (Mux29)))) # (!Selector5 & (((\Selector61~0_combout ))))

	.dataa(\rf|Mux29~20_combout ),
	.datab(\cu|Selector5~2_combout ),
	.datac(dcifimemload_0),
	.datad(\Selector61~0_combout ),
	.cin(gnd),
	.combout(\Selector61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector61~1 .lut_mask = 16'hF388;
defparam \Selector61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N10
cycloneive_lcell_comb \Selector58~0 (
// Equation(s):
// \Selector58~0_combout  = (Selector5 & (((Selector6) # (Mux26)))) # (!Selector5 & (\Add1~6_combout  & (!Selector6)))

	.dataa(\Add1~6_combout ),
	.datab(\cu|Selector5~2_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\rf|Mux26~20_combout ),
	.cin(gnd),
	.combout(\Selector58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector58~0 .lut_mask = 16'hCEC2;
defparam \Selector58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N0
cycloneive_lcell_comb \Selector58~1 (
// Equation(s):
// \Selector58~1_combout  = (Selector6 & ((\Selector58~0_combout  & (dcifimemload_3)) # (!\Selector58~0_combout  & ((\Add2~6_combout ))))) # (!Selector6 & (((\Selector58~0_combout ))))

	.dataa(dcifimemload_3),
	.datab(\Add2~6_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Selector58~0_combout ),
	.cin(gnd),
	.combout(\Selector58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector58~1 .lut_mask = 16'hAFC0;
defparam \Selector58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N10
cycloneive_lcell_comb \Selector59~0 (
// Equation(s):
// \Selector59~0_combout  = (Selector6 & (((\Add2~4_combout ) # (Selector5)))) # (!Selector6 & (\Add1~4_combout  & ((!Selector5))))

	.dataa(\Add1~4_combout ),
	.datab(\Add2~4_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\cu|Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector59~0 .lut_mask = 16'hF0CA;
defparam \Selector59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N28
cycloneive_lcell_comb \Selector59~1 (
// Equation(s):
// \Selector59~1_combout  = (Selector5 & ((\Selector59~0_combout  & (dcifimemload_2)) # (!\Selector59~0_combout  & ((Mux27))))) # (!Selector5 & (((\Selector59~0_combout ))))

	.dataa(dcifimemload_2),
	.datab(\rf|Mux27~20_combout ),
	.datac(\cu|Selector5~2_combout ),
	.datad(\Selector59~0_combout ),
	.cin(gnd),
	.combout(\Selector59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector59~1 .lut_mask = 16'hAFC0;
defparam \Selector59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N20
cycloneive_lcell_comb \Selector56~0 (
// Equation(s):
// \Selector56~0_combout  = (Selector6 & (((Selector5)))) # (!Selector6 & ((Selector5 & ((Mux24))) # (!Selector5 & (\Add1~10_combout ))))

	.dataa(\Add1~10_combout ),
	.datab(\rf|Mux24~20_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\cu|Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector56~0 .lut_mask = 16'hFC0A;
defparam \Selector56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N4
cycloneive_lcell_comb \Selector56~1 (
// Equation(s):
// \Selector56~1_combout  = (Selector6 & ((\Selector56~0_combout  & ((dcifimemload_5))) # (!\Selector56~0_combout  & (\Add2~10_combout )))) # (!Selector6 & (((\Selector56~0_combout ))))

	.dataa(\cu|Selector6~1_combout ),
	.datab(\Add2~10_combout ),
	.datac(dcifimemload_5),
	.datad(\Selector56~0_combout ),
	.cin(gnd),
	.combout(\Selector56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector56~1 .lut_mask = 16'hF588;
defparam \Selector56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N22
cycloneive_lcell_comb \Selector57~0 (
// Equation(s):
// \Selector57~0_combout  = (Selector6 & ((\Add2~8_combout ) # ((Selector5)))) # (!Selector6 & (((\Add1~8_combout  & !Selector5))))

	.dataa(\Add2~8_combout ),
	.datab(\Add1~8_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\cu|Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector57~0 .lut_mask = 16'hF0AC;
defparam \Selector57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N6
cycloneive_lcell_comb \Selector57~1 (
// Equation(s):
// \Selector57~1_combout  = (\Selector57~0_combout  & (((dcifimemload_4) # (!Selector5)))) # (!\Selector57~0_combout  & (Mux25 & ((Selector5))))

	.dataa(\rf|Mux25~20_combout ),
	.datab(dcifimemload_4),
	.datac(\Selector57~0_combout ),
	.datad(\cu|Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector57~1 .lut_mask = 16'hCAF0;
defparam \Selector57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N10
cycloneive_lcell_comb \Selector54~0 (
// Equation(s):
// \Selector54~0_combout  = (Selector5 & (((Mux22) # (Selector6)))) # (!Selector5 & (\Add1~14_combout  & ((!Selector6))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\Add1~14_combout ),
	.datac(\rf|Mux22~20_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector54~0 .lut_mask = 16'hAAE4;
defparam \Selector54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N26
cycloneive_lcell_comb \Selector54~1 (
// Equation(s):
// \Selector54~1_combout  = (Selector6 & ((\Selector54~0_combout  & ((dcifimemload_7))) # (!\Selector54~0_combout  & (\Add2~14_combout )))) # (!Selector6 & (((\Selector54~0_combout ))))

	.dataa(\Add2~14_combout ),
	.datab(dcifimemload_7),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Selector54~0_combout ),
	.cin(gnd),
	.combout(\Selector54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector54~1 .lut_mask = 16'hCFA0;
defparam \Selector54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N20
cycloneive_lcell_comb \Selector55~0 (
// Equation(s):
// \Selector55~0_combout  = (Selector6 & (((\Add2~12_combout ) # (Selector5)))) # (!Selector6 & (\Add1~12_combout  & ((!Selector5))))

	.dataa(\Add1~12_combout ),
	.datab(\Add2~12_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\cu|Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector55~0 .lut_mask = 16'hF0CA;
defparam \Selector55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N8
cycloneive_lcell_comb \Selector55~1 (
// Equation(s):
// \Selector55~1_combout  = (Selector5 & ((\Selector55~0_combout  & (dcifimemload_6)) # (!\Selector55~0_combout  & ((Mux23))))) # (!Selector5 & (((\Selector55~0_combout ))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(dcifimemload_6),
	.datac(\rf|Mux23~20_combout ),
	.datad(\Selector55~0_combout ),
	.cin(gnd),
	.combout(\Selector55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector55~1 .lut_mask = 16'hDDA0;
defparam \Selector55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N6
cycloneive_lcell_comb \Selector52~0 (
// Equation(s):
// \Selector52~0_combout  = (Selector5 & (((Mux20) # (Selector6)))) # (!Selector5 & (\Add1~18_combout  & ((!Selector6))))

	.dataa(\Add1~18_combout ),
	.datab(\rf|Mux20~20_combout ),
	.datac(\cu|Selector5~2_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector52~0 .lut_mask = 16'hF0CA;
defparam \Selector52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N24
cycloneive_lcell_comb \Selector52~1 (
// Equation(s):
// \Selector52~1_combout  = (Selector6 & ((\Selector52~0_combout  & ((dcifimemload_9))) # (!\Selector52~0_combout  & (\Add2~18_combout )))) # (!Selector6 & (((\Selector52~0_combout ))))

	.dataa(\Add2~18_combout ),
	.datab(\cu|Selector6~1_combout ),
	.datac(dcifimemload_9),
	.datad(\Selector52~0_combout ),
	.cin(gnd),
	.combout(\Selector52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector52~1 .lut_mask = 16'hF388;
defparam \Selector52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N16
cycloneive_lcell_comb \Selector53~0 (
// Equation(s):
// \Selector53~0_combout  = (Selector5 & (((Selector6)))) # (!Selector5 & ((Selector6 & (\Add2~16_combout )) # (!Selector6 & ((\Add1~16_combout )))))

	.dataa(\Add2~16_combout ),
	.datab(\Add1~16_combout ),
	.datac(\cu|Selector5~2_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector53~0 .lut_mask = 16'hFA0C;
defparam \Selector53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N26
cycloneive_lcell_comb \Selector53~1 (
// Equation(s):
// \Selector53~1_combout  = (Selector5 & ((\Selector53~0_combout  & (dcifimemload_8)) # (!\Selector53~0_combout  & ((Mux21))))) # (!Selector5 & (((\Selector53~0_combout ))))

	.dataa(dcifimemload_8),
	.datab(\rf|Mux21~20_combout ),
	.datac(\cu|Selector5~2_combout ),
	.datad(\Selector53~0_combout ),
	.cin(gnd),
	.combout(\Selector53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector53~1 .lut_mask = 16'hAFC0;
defparam \Selector53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N28
cycloneive_lcell_comb \Selector50~0 (
// Equation(s):
// \Selector50~0_combout  = (Selector5 & ((Mux18) # ((Selector6)))) # (!Selector5 & (((\Add1~22_combout  & !Selector6))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\rf|Mux18~20_combout ),
	.datac(\Add1~22_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector50~0 .lut_mask = 16'hAAD8;
defparam \Selector50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N8
cycloneive_lcell_comb \Selector50~1 (
// Equation(s):
// \Selector50~1_combout  = (Selector6 & ((\Selector50~0_combout  & (dcifimemload_11)) # (!\Selector50~0_combout  & ((\Add2~22_combout ))))) # (!Selector6 & (((\Selector50~0_combout ))))

	.dataa(dcifimemload_11),
	.datab(\Add2~22_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Selector50~0_combout ),
	.cin(gnd),
	.combout(\Selector50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector50~1 .lut_mask = 16'hAFC0;
defparam \Selector50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N10
cycloneive_lcell_comb \Selector51~0 (
// Equation(s):
// \Selector51~0_combout  = (Selector5 & (((Selector6)))) # (!Selector5 & ((Selector6 & (\Add2~20_combout )) # (!Selector6 & ((\Add1~20_combout )))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\Add2~20_combout ),
	.datac(\Add1~20_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector51~0 .lut_mask = 16'hEE50;
defparam \Selector51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N30
cycloneive_lcell_comb \Selector51~1 (
// Equation(s):
// \Selector51~1_combout  = (Selector5 & ((\Selector51~0_combout  & (dcifimemload_10)) # (!\Selector51~0_combout  & ((Mux19))))) # (!Selector5 & (((\Selector51~0_combout ))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(dcifimemload_10),
	.datac(\rf|Mux19~20_combout ),
	.datad(\Selector51~0_combout ),
	.cin(gnd),
	.combout(\Selector51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector51~1 .lut_mask = 16'hDDA0;
defparam \Selector51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N4
cycloneive_lcell_comb \Selector48~0 (
// Equation(s):
// \Selector48~0_combout  = (Selector5 & (((Mux16) # (Selector6)))) # (!Selector5 & (\Add1~26_combout  & ((!Selector6))))

	.dataa(\Add1~26_combout ),
	.datab(\rf|Mux16~20_combout ),
	.datac(\cu|Selector5~2_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector48~0 .lut_mask = 16'hF0CA;
defparam \Selector48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N12
cycloneive_lcell_comb \Selector48~1 (
// Equation(s):
// \Selector48~1_combout  = (\Selector48~0_combout  & ((dcifimemload_13) # ((!Selector6)))) # (!\Selector48~0_combout  & (((\Add2~26_combout  & Selector6))))

	.dataa(dcifimemload_13),
	.datab(\Add2~26_combout ),
	.datac(\Selector48~0_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector48~1 .lut_mask = 16'hACF0;
defparam \Selector48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N18
cycloneive_lcell_comb \Selector49~0 (
// Equation(s):
// \Selector49~0_combout  = (Selector5 & (((Selector6)))) # (!Selector5 & ((Selector6 & (\Add2~24_combout )) # (!Selector6 & ((\Add1~24_combout )))))

	.dataa(\Add2~24_combout ),
	.datab(\Add1~24_combout ),
	.datac(\cu|Selector5~2_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector49~0 .lut_mask = 16'hFA0C;
defparam \Selector49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N22
cycloneive_lcell_comb \Selector49~1 (
// Equation(s):
// \Selector49~1_combout  = (Selector5 & ((\Selector49~0_combout  & (dcifimemload_12)) # (!\Selector49~0_combout  & ((Mux17))))) # (!Selector5 & (((\Selector49~0_combout ))))

	.dataa(dcifimemload_12),
	.datab(\rf|Mux17~20_combout ),
	.datac(\cu|Selector5~2_combout ),
	.datad(\Selector49~0_combout ),
	.cin(gnd),
	.combout(\Selector49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector49~1 .lut_mask = 16'hAFC0;
defparam \Selector49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N4
cycloneive_lcell_comb \Selector46~0 (
// Equation(s):
// \Selector46~0_combout  = (Selector5 & ((Selector6) # ((Mux14)))) # (!Selector5 & (!Selector6 & (\Add1~30_combout )))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\cu|Selector6~1_combout ),
	.datac(\Add1~30_combout ),
	.datad(\rf|Mux14~20_combout ),
	.cin(gnd),
	.combout(\Selector46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector46~0 .lut_mask = 16'hBA98;
defparam \Selector46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N20
cycloneive_lcell_comb \Selector46~1 (
// Equation(s):
// \Selector46~1_combout  = (Selector6 & ((\Selector46~0_combout  & ((dcifimemload_15))) # (!\Selector46~0_combout  & (\Add2~30_combout )))) # (!Selector6 & (((\Selector46~0_combout ))))

	.dataa(\Add2~30_combout ),
	.datab(\cu|Selector6~1_combout ),
	.datac(\Selector46~0_combout ),
	.datad(dcifimemload_15),
	.cin(gnd),
	.combout(\Selector46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector46~1 .lut_mask = 16'hF838;
defparam \Selector46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N10
cycloneive_lcell_comb \Selector47~0 (
// Equation(s):
// \Selector47~0_combout  = (Selector5 & (((Selector6)))) # (!Selector5 & ((Selector6 & ((\Add2~28_combout ))) # (!Selector6 & (\Add1~28_combout ))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\Add1~28_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Add2~28_combout ),
	.cin(gnd),
	.combout(\Selector47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector47~0 .lut_mask = 16'hF4A4;
defparam \Selector47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N30
cycloneive_lcell_comb \Selector47~1 (
// Equation(s):
// \Selector47~1_combout  = (Selector5 & ((\Selector47~0_combout  & ((dcifimemload_14))) # (!\Selector47~0_combout  & (Mux15)))) # (!Selector5 & (((\Selector47~0_combout ))))

	.dataa(\rf|Mux15~20_combout ),
	.datab(dcifimemload_14),
	.datac(\cu|Selector5~2_combout ),
	.datad(\Selector47~0_combout ),
	.cin(gnd),
	.combout(\Selector47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector47~1 .lut_mask = 16'hCFA0;
defparam \Selector47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N28
cycloneive_lcell_comb \Selector44~0 (
// Equation(s):
// \Selector44~0_combout  = (Selector6 & (((Selector5)))) # (!Selector6 & ((Selector5 & (Mux12)) # (!Selector5 & ((\Add1~34_combout )))))

	.dataa(\rf|Mux12~20_combout ),
	.datab(\Add1~34_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\cu|Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector44~0 .lut_mask = 16'hFA0C;
defparam \Selector44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N4
cycloneive_lcell_comb \Selector44~1 (
// Equation(s):
// \Selector44~1_combout  = (Selector6 & ((\Selector44~0_combout  & ((dcifimemload_17))) # (!\Selector44~0_combout  & (\Add2~34_combout )))) # (!Selector6 & (((\Selector44~0_combout ))))

	.dataa(\cu|Selector6~1_combout ),
	.datab(\Add2~34_combout ),
	.datac(dcifimemload_17),
	.datad(\Selector44~0_combout ),
	.cin(gnd),
	.combout(\Selector44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector44~1 .lut_mask = 16'hF588;
defparam \Selector44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N14
cycloneive_lcell_comb \Selector45~0 (
// Equation(s):
// \Selector45~0_combout  = (Selector6 & ((\Add2~32_combout ) # ((Selector5)))) # (!Selector6 & (((\Add1~32_combout  & !Selector5))))

	.dataa(\Add2~32_combout ),
	.datab(\Add1~32_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\cu|Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector45~0 .lut_mask = 16'hF0AC;
defparam \Selector45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N12
cycloneive_lcell_comb \Selector45~1 (
// Equation(s):
// \Selector45~1_combout  = (Selector5 & ((\Selector45~0_combout  & (dcifimemload_16)) # (!\Selector45~0_combout  & ((Mux13))))) # (!Selector5 & (((\Selector45~0_combout ))))

	.dataa(dcifimemload_16),
	.datab(\cu|Selector5~2_combout ),
	.datac(\Selector45~0_combout ),
	.datad(\rf|Mux13~20_combout ),
	.cin(gnd),
	.combout(\Selector45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector45~1 .lut_mask = 16'hBCB0;
defparam \Selector45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N10
cycloneive_lcell_comb \Selector42~0 (
// Equation(s):
// \Selector42~0_combout  = (Selector5 & ((Mux10) # ((Selector6)))) # (!Selector5 & (((!Selector6 & \Add1~38_combout ))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\rf|Mux10~20_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Add1~38_combout ),
	.cin(gnd),
	.combout(\Selector42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector42~0 .lut_mask = 16'hADA8;
defparam \Selector42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N4
cycloneive_lcell_comb \Selector42~1 (
// Equation(s):
// \Selector42~1_combout  = (Selector6 & ((\Selector42~0_combout  & (dcifimemload_19)) # (!\Selector42~0_combout  & ((\Add2~38_combout ))))) # (!Selector6 & (((\Selector42~0_combout ))))

	.dataa(\cu|Selector6~1_combout ),
	.datab(dcifimemload_19),
	.datac(\Add2~38_combout ),
	.datad(\Selector42~0_combout ),
	.cin(gnd),
	.combout(\Selector42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector42~1 .lut_mask = 16'hDDA0;
defparam \Selector42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N12
cycloneive_lcell_comb \Selector43~0 (
// Equation(s):
// \Selector43~0_combout  = (Selector5 & (((Selector6)))) # (!Selector5 & ((Selector6 & ((\Add2~36_combout ))) # (!Selector6 & (\Add1~36_combout ))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\Add1~36_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Add2~36_combout ),
	.cin(gnd),
	.combout(\Selector43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector43~0 .lut_mask = 16'hF4A4;
defparam \Selector43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N26
cycloneive_lcell_comb \Selector43~1 (
// Equation(s):
// \Selector43~1_combout  = (Selector5 & ((\Selector43~0_combout  & ((dcifimemload_18))) # (!\Selector43~0_combout  & (Mux11)))) # (!Selector5 & (((\Selector43~0_combout ))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\rf|Mux11~20_combout ),
	.datac(dcifimemload_18),
	.datad(\Selector43~0_combout ),
	.cin(gnd),
	.combout(\Selector43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector43~1 .lut_mask = 16'hF588;
defparam \Selector43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N8
cycloneive_lcell_comb \Selector40~0 (
// Equation(s):
// \Selector40~0_combout  = (Selector5 & ((Mux8) # ((Selector6)))) # (!Selector5 & (((\Add1~42_combout  & !Selector6))))

	.dataa(\rf|Mux8~20_combout ),
	.datab(\cu|Selector5~2_combout ),
	.datac(\Add1~42_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector40~0 .lut_mask = 16'hCCB8;
defparam \Selector40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N4
cycloneive_lcell_comb \Selector40~1 (
// Equation(s):
// \Selector40~1_combout  = (\Selector40~0_combout  & (((dcifimemload_21) # (!Selector6)))) # (!\Selector40~0_combout  & (\Add2~42_combout  & ((Selector6))))

	.dataa(\Add2~42_combout ),
	.datab(dcifimemload_21),
	.datac(\Selector40~0_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector40~1 .lut_mask = 16'hCAF0;
defparam \Selector40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N2
cycloneive_lcell_comb \Selector41~0 (
// Equation(s):
// \Selector41~0_combout  = (Selector5 & (((Selector6)))) # (!Selector5 & ((Selector6 & (\Add2~40_combout )) # (!Selector6 & ((\Add1~40_combout )))))

	.dataa(\Add2~40_combout ),
	.datab(\Add1~40_combout ),
	.datac(\cu|Selector5~2_combout ),
	.datad(\cu|Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector41~0 .lut_mask = 16'hFA0C;
defparam \Selector41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N30
cycloneive_lcell_comb \Selector41~1 (
// Equation(s):
// \Selector41~1_combout  = (Selector5 & ((\Selector41~0_combout  & ((dcifimemload_20))) # (!\Selector41~0_combout  & (Mux9)))) # (!Selector5 & (((\Selector41~0_combout ))))

	.dataa(\rf|Mux9~20_combout ),
	.datab(\cu|Selector5~2_combout ),
	.datac(dcifimemload_20),
	.datad(\Selector41~0_combout ),
	.cin(gnd),
	.combout(\Selector41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector41~1 .lut_mask = 16'hF388;
defparam \Selector41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N12
cycloneive_lcell_comb \Selector38~0 (
// Equation(s):
// \Selector38~0_combout  = (Selector5 & ((Mux6) # ((Selector6)))) # (!Selector5 & (((!Selector6 & \Add1~46_combout ))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(\rf|Mux6~20_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Add1~46_combout ),
	.cin(gnd),
	.combout(\Selector38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector38~0 .lut_mask = 16'hADA8;
defparam \Selector38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N4
cycloneive_lcell_comb \Selector38~1 (
// Equation(s):
// \Selector38~1_combout  = (Selector6 & ((\Selector38~0_combout  & (dcifimemload_23)) # (!\Selector38~0_combout  & ((\Add2~46_combout ))))) # (!Selector6 & (((\Selector38~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Add2~46_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Selector38~0_combout ),
	.cin(gnd),
	.combout(\Selector38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector38~1 .lut_mask = 16'hAFC0;
defparam \Selector38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N10
cycloneive_lcell_comb \Selector39~0 (
// Equation(s):
// \Selector39~0_combout  = (Selector5 & (((Selector6)))) # (!Selector5 & ((Selector6 & ((\Add2~44_combout ))) # (!Selector6 & (\Add1~44_combout ))))

	.dataa(\Add1~44_combout ),
	.datab(\cu|Selector5~2_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Add2~44_combout ),
	.cin(gnd),
	.combout(\Selector39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector39~0 .lut_mask = 16'hF2C2;
defparam \Selector39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N26
cycloneive_lcell_comb \Selector39~1 (
// Equation(s):
// \Selector39~1_combout  = (Selector5 & ((\Selector39~0_combout  & (dcifimemload_22)) # (!\Selector39~0_combout  & ((Mux7))))) # (!Selector5 & (((\Selector39~0_combout ))))

	.dataa(\cu|Selector5~2_combout ),
	.datab(dcifimemload_22),
	.datac(\rf|Mux7~20_combout ),
	.datad(\Selector39~0_combout ),
	.cin(gnd),
	.combout(\Selector39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector39~1 .lut_mask = 16'hDDA0;
defparam \Selector39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N12
cycloneive_lcell_comb \Selector36~0 (
// Equation(s):
// \Selector36~0_combout  = (Selector6 & (((Selector5)))) # (!Selector6 & ((Selector5 & ((Mux4))) # (!Selector5 & (\Add1~50_combout ))))

	.dataa(\Add1~50_combout ),
	.datab(\rf|Mux4~20_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\cu|Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector36~0 .lut_mask = 16'hFC0A;
defparam \Selector36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N26
cycloneive_lcell_comb \Selector36~1 (
// Equation(s):
// \Selector36~1_combout  = (Selector6 & ((\Selector36~0_combout  & (dcifimemload_25)) # (!\Selector36~0_combout  & ((\Add2~50_combout ))))) # (!Selector6 & (((\Selector36~0_combout ))))

	.dataa(dcifimemload_25),
	.datab(\Add2~50_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Selector36~0_combout ),
	.cin(gnd),
	.combout(\Selector36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector36~1 .lut_mask = 16'hAFC0;
defparam \Selector36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N6
cycloneive_lcell_comb \Selector37~0 (
// Equation(s):
// \Selector37~0_combout  = (Selector5 & (((Selector6)))) # (!Selector5 & ((Selector6 & ((\Add2~48_combout ))) # (!Selector6 & (\Add1~48_combout ))))

	.dataa(\Add1~48_combout ),
	.datab(\cu|Selector5~2_combout ),
	.datac(\cu|Selector6~1_combout ),
	.datad(\Add2~48_combout ),
	.cin(gnd),
	.combout(\Selector37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector37~0 .lut_mask = 16'hF2C2;
defparam \Selector37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N4
cycloneive_lcell_comb \Selector37~1 (
// Equation(s):
// \Selector37~1_combout  = (Selector5 & ((\Selector37~0_combout  & ((dcifimemload_24))) # (!\Selector37~0_combout  & (Mux5)))) # (!Selector5 & (((\Selector37~0_combout ))))

	.dataa(\rf|Mux5~20_combout ),
	.datab(\cu|Selector5~2_combout ),
	.datac(dcifimemload_24),
	.datad(\Selector37~0_combout ),
	.cin(gnd),
	.combout(\Selector37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector37~1 .lut_mask = 16'hF388;
defparam \Selector37~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu (
	Mux63,
	Mux30,
	Selector95,
	Mux33,
	Selector70,
	Selector3,
	Mux1,
	Mux34,
	Selector71,
	Mux2,
	Mux35,
	Selector72,
	Mux3,
	Mux36,
	Selector73,
	Mux4,
	Mux37,
	Selector74,
	Mux5,
	Mux38,
	Selector75,
	Mux6,
	Mux39,
	Selector76,
	Mux7,
	Mux40,
	Selector77,
	Mux8,
	Mux41,
	Selector78,
	Mux9,
	Mux42,
	Selector79,
	Mux10,
	Mux43,
	Selector80,
	Mux11,
	Mux44,
	Selector81,
	Mux12,
	Mux45,
	Selector82,
	Mux13,
	Mux46,
	Selector83,
	Mux14,
	Mux47,
	Selector84,
	Mux15,
	Mux48,
	Selector85,
	Mux16,
	Mux49,
	Selector86,
	Mux17,
	Mux50,
	Selector87,
	Mux18,
	Mux51,
	Selector88,
	Mux19,
	Mux52,
	Selector89,
	Mux20,
	Mux53,
	Selector90,
	Mux21,
	Mux54,
	Selector91,
	Mux22,
	Mux55,
	Selector92,
	Mux23,
	Mux56,
	Selector93,
	Mux24,
	Mux57,
	Selector94,
	Mux25,
	Mux58,
	Selector951,
	Mux26,
	Selector100,
	Mux59,
	Selector96,
	Mux27,
	Mux60,
	Selector97,
	Mux28,
	Mux61,
	Selector98,
	Mux29,
	Mux62,
	Selector99,
	Selector1001,
	Mux31,
	Selector991,
	Selector1002,
	Selector981,
	Selector952,
	Selector941,
	Selector931,
	Selector921,
	Selector911,
	Selector901,
	Selector891,
	Selector881,
	Selector871,
	Selector861,
	Selector851,
	Selector841,
	Selector831,
	Selector821,
	Selector811,
	Selector801,
	Selector791,
	Selector781,
	Selector771,
	Selector761,
	Selector751,
	Selector741,
	Selector731,
	Selector721,
	Selector711,
	Selector701,
	Selector69,
	Mux32,
	Selector691,
	Selector961,
	Mux0,
	Selector971,
	Selector0,
	Selector1,
	Selector2,
	Mux110,
	Mux311,
	Mux111,
	Mux01,
	Mux02,
	Mux241,
	Mux251,
	Mux261,
	Mux271,
	Mux410,
	Mux510,
	Mux64,
	Mux71,
	Equal0,
	Mux310,
	Mux210,
	Mux231,
	Mux232,
	Mux221,
	Mux222,
	Mux211,
	Mux212,
	Mux201,
	Mux202,
	Mux191,
	Mux192,
	Mux181,
	Mux182,
	Mux171,
	Mux172,
	Mux161,
	Mux162,
	Mux291,
	Mux281,
	Mux81,
	Mux101,
	Mux102,
	Mux91,
	Mux92,
	Mux301,
	Mux151,
	Mux152,
	Mux141,
	Mux142,
	Mux131,
	Mux132,
	Mux121,
	Mux122,
	Mux112,
	Mux113,
	Equal01,
	Mux312,
	Mux114,
	Mux03,
	Mux233,
	Mux223,
	Mux213,
	Mux203,
	Mux193,
	Mux183,
	Mux173,
	Mux163,
	Mux103,
	Mux93,
	Mux153,
	Mux143,
	Mux133,
	Mux123,
	Mux115,
	devpor,
	devclrn,
	devoe);
input 	Mux63;
input 	Mux30;
input 	Selector95;
input 	Mux33;
input 	Selector70;
input 	Selector3;
input 	Mux1;
input 	Mux34;
input 	Selector71;
input 	Mux2;
input 	Mux35;
input 	Selector72;
input 	Mux3;
input 	Mux36;
input 	Selector73;
input 	Mux4;
input 	Mux37;
input 	Selector74;
input 	Mux5;
input 	Mux38;
input 	Selector75;
input 	Mux6;
input 	Mux39;
input 	Selector76;
input 	Mux7;
input 	Mux40;
input 	Selector77;
input 	Mux8;
input 	Mux41;
input 	Selector78;
input 	Mux9;
input 	Mux42;
input 	Selector79;
input 	Mux10;
input 	Mux43;
input 	Selector80;
input 	Mux11;
input 	Mux44;
input 	Selector81;
input 	Mux12;
input 	Mux45;
input 	Selector82;
input 	Mux13;
input 	Mux46;
input 	Selector83;
input 	Mux14;
input 	Mux47;
input 	Selector84;
input 	Mux15;
input 	Mux48;
input 	Selector85;
input 	Mux16;
input 	Mux49;
input 	Selector86;
input 	Mux17;
input 	Mux50;
input 	Selector87;
input 	Mux18;
input 	Mux51;
input 	Selector88;
input 	Mux19;
input 	Mux52;
input 	Selector89;
input 	Mux20;
input 	Mux53;
input 	Selector90;
input 	Mux21;
input 	Mux54;
input 	Selector91;
input 	Mux22;
input 	Mux55;
input 	Selector92;
input 	Mux23;
input 	Mux56;
input 	Selector93;
input 	Mux24;
input 	Mux57;
input 	Selector94;
input 	Mux25;
input 	Mux58;
input 	Selector951;
input 	Mux26;
input 	Selector100;
input 	Mux59;
input 	Selector96;
input 	Mux27;
input 	Mux60;
input 	Selector97;
input 	Mux28;
input 	Mux61;
input 	Selector98;
input 	Mux29;
input 	Mux62;
input 	Selector99;
input 	Selector1001;
input 	Mux31;
input 	Selector991;
input 	Selector1002;
input 	Selector981;
input 	Selector952;
input 	Selector941;
input 	Selector931;
input 	Selector921;
input 	Selector911;
input 	Selector901;
input 	Selector891;
input 	Selector881;
input 	Selector871;
input 	Selector861;
input 	Selector851;
input 	Selector841;
input 	Selector831;
input 	Selector821;
input 	Selector811;
input 	Selector801;
input 	Selector791;
input 	Selector781;
input 	Selector771;
input 	Selector761;
input 	Selector751;
input 	Selector741;
input 	Selector731;
input 	Selector721;
input 	Selector711;
input 	Selector701;
input 	Selector69;
input 	Mux32;
input 	Selector691;
input 	Selector961;
input 	Mux0;
input 	Selector971;
input 	Selector0;
input 	Selector1;
input 	Selector2;
output 	Mux110;
output 	Mux311;
output 	Mux111;
output 	Mux01;
output 	Mux02;
output 	Mux241;
output 	Mux251;
output 	Mux261;
output 	Mux271;
output 	Mux410;
output 	Mux510;
output 	Mux64;
output 	Mux71;
output 	Equal0;
output 	Mux310;
output 	Mux210;
output 	Mux231;
output 	Mux232;
output 	Mux221;
output 	Mux222;
output 	Mux211;
output 	Mux212;
output 	Mux201;
output 	Mux202;
output 	Mux191;
output 	Mux192;
output 	Mux181;
output 	Mux182;
output 	Mux171;
output 	Mux172;
output 	Mux161;
output 	Mux162;
output 	Mux291;
output 	Mux281;
output 	Mux81;
output 	Mux101;
output 	Mux102;
output 	Mux91;
output 	Mux92;
output 	Mux301;
output 	Mux151;
output 	Mux152;
output 	Mux141;
output 	Mux142;
output 	Mux131;
output 	Mux132;
output 	Mux121;
output 	Mux122;
output 	Mux112;
output 	Mux113;
output 	Equal01;
output 	Mux312;
output 	Mux114;
output 	Mux03;
output 	Mux233;
output 	Mux223;
output 	Mux213;
output 	Mux203;
output 	Mux193;
output 	Mux183;
output 	Mux173;
output 	Mux163;
output 	Mux103;
output 	Mux93;
output 	Mux153;
output 	Mux143;
output 	Mux133;
output 	Mux123;
output 	Mux115;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add0~37_combout ;
wire \Add0~39_combout ;
wire \Add0~1_combout ;
wire \Add0~2_combout ;
wire \Add0~3_combout ;
wire \Add0~5_combout ;
wire \Add0~7_combout ;
wire \Add0~25_combout ;
wire \Add0~26_combout ;
wire \Add0~27_combout ;
wire \Add0~28_combout ;
wire \Add0~29_combout ;
wire \Add0~30_combout ;
wire \ShiftLeft0~11_combout ;
wire \ShiftRight0~37_combout ;
wire \ShiftRight0~38_combout ;
wire \ShiftLeft0~80_combout ;
wire \Mux2~6_combout ;
wire \Mux19~2_combout ;
wire \Mux18~5_combout ;
wire \Mux15~3_combout ;
wire \Mux11~2_combout ;
wire \Mux8~10_combout ;
wire \Mux9~8_combout ;
wire \Mux23~3_combout ;
wire \Mux23~2_combout ;
wire \ShiftLeft0~17_combout ;
wire \ShiftLeft0~18_combout ;
wire \ShiftLeft0~16_combout ;
wire \ShiftLeft0~12_combout ;
wire \ShiftLeft0~14_combout ;
wire \ShiftLeft0~13_combout ;
wire \ShiftLeft0~15_combout ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \ShiftLeft0~4_combout ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~5_combout ;
wire \ShiftLeft0~1_combout ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~2_combout ;
wire \ShiftLeft0~6_combout ;
wire \Mux0~2_combout ;
wire \ShiftLeft0~8_combout ;
wire \ShiftLeft0~9_combout ;
wire \ShiftLeft0~10_combout ;
wire \ShiftLeft0~7_combout ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux0~6_combout ;
wire \ShiftLeft0~22_combout ;
wire \ShiftLeft0~23_combout ;
wire \ShiftLeft0~19_combout ;
wire \ShiftLeft0~20_combout ;
wire \ShiftLeft0~24_combout ;
wire \ShiftLeft0~29_combout ;
wire \ShiftLeft0~30_combout ;
wire \ShiftLeft0~25_combout ;
wire \ShiftLeft0~26_combout ;
wire \ShiftLeft0~27_combout ;
wire \ShiftLeft0~31_combout ;
wire \ShiftLeft0~32_combout ;
wire \Mux1~4_combout ;
wire \ShiftRight0~6_combout ;
wire \ShiftRight0~103_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \Add0~0_combout ;
wire \Add0~4_combout ;
wire \Add0~6_combout ;
wire \Add0~13_combout ;
wire \Add0~15_combout ;
wire \Add0~16_combout ;
wire \Add0~17_combout ;
wire \Add0~19_combout ;
wire \Add0~20_combout ;
wire \Add0~23_combout ;
wire \Add0~24_combout ;
wire \Add0~32_cout ;
wire \Add0~34 ;
wire \Add0~36 ;
wire \Add0~38 ;
wire \Add0~40 ;
wire \Add0~42 ;
wire \Add0~44 ;
wire \Add0~46 ;
wire \Add0~48 ;
wire \Add0~50 ;
wire \Add0~52 ;
wire \Add0~54 ;
wire \Add0~56 ;
wire \Add0~58 ;
wire \Add0~60 ;
wire \Add0~62 ;
wire \Add0~64 ;
wire \Add0~66 ;
wire \Add0~68 ;
wire \Add0~70 ;
wire \Add0~72 ;
wire \Add0~74 ;
wire \Add0~76 ;
wire \Add0~78 ;
wire \Add0~80 ;
wire \Add0~82 ;
wire \Add0~84 ;
wire \Add0~86 ;
wire \Add0~88 ;
wire \Add0~90 ;
wire \Add0~92 ;
wire \Add0~93_combout ;
wire \Mux0~3_combout ;
wire \ShiftLeft0~38_combout ;
wire \Mux0~8_combout ;
wire \Mux0~9_combout ;
wire \ShiftLeft0~35_combout ;
wire \ShiftLeft0~36_combout ;
wire \ShiftLeft0~33_combout ;
wire \ShiftLeft0~34_combout ;
wire \ShiftLeft0~37_combout ;
wire \ShiftRight0~7_combout ;
wire \ShiftLeft0~42_combout ;
wire \ShiftLeft0~43_combout ;
wire \ShiftLeft0~44_combout ;
wire \ShiftLeft0~45_combout ;
wire \ShiftLeft0~46_combout ;
wire \ShiftLeft0~47_combout ;
wire \ShiftLeft0~48_combout ;
wire \ShiftLeft0~49_combout ;
wire \ShiftLeft0~50_combout ;
wire \ShiftLeft0~51_combout ;
wire \ShiftLeft0~52_combout ;
wire \Mux0~10_combout ;
wire \Mux0~11_combout ;
wire \Mux0~12_combout ;
wire \Add0~95_combout ;
wire \Add0~94 ;
wire \Add0~96_combout ;
wire \Mux24~10_combout ;
wire \Mux24~7_combout ;
wire \Mux30~0_combout ;
wire \Mux6~11_combout ;
wire \Add0~47_combout ;
wire \Mux24~8_combout ;
wire \Mux24~6_combout ;
wire \Mux6~18_combout ;
wire \ShiftRight0~16_combout ;
wire \ShiftRight0~15_combout ;
wire \ShiftRight0~17_combout ;
wire \Mux6~10_combout ;
wire \Mux24~4_combout ;
wire \ShiftRight0~12_combout ;
wire \ShiftRight0~11_combout ;
wire \ShiftRight0~13_combout ;
wire \ShiftRight0~8_combout ;
wire \ShiftRight0~9_combout ;
wire \ShiftRight0~10_combout ;
wire \ShiftRight0~14_combout ;
wire \ShiftRight0~21_combout ;
wire \ShiftRight0~22_combout ;
wire \ShiftRight0~23_combout ;
wire \ShiftRight0~24_combout ;
wire \ShiftRight0~25_combout ;
wire \ShiftRight0~26_combout ;
wire \ShiftRight0~27_combout ;
wire \ShiftRight0~28_combout ;
wire \ShiftRight0~29_combout ;
wire \Mux24~5_combout ;
wire \Mux25~2_combout ;
wire \ShiftRight0~39_combout ;
wire \ShiftRight0~40_combout ;
wire \ShiftRight0~41_combout ;
wire \ShiftRight0~42_combout ;
wire \ShiftRight0~43_combout ;
wire \ShiftRight0~44_combout ;
wire \ShiftRight0~30_combout ;
wire \ShiftRight0~31_combout ;
wire \ShiftRight0~32_combout ;
wire \ShiftRight0~33_combout ;
wire \ShiftRight0~34_combout ;
wire \ShiftRight0~35_combout ;
wire \ShiftRight0~36_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux25~3_combout ;
wire \Add0~45_combout ;
wire \Mux25~4_combout ;
wire \Mux26~3_combout ;
wire \Add0~43_combout ;
wire \Mux26~4_combout ;
wire \ShiftLeft0~53_combout ;
wire \ShiftLeft0~21_combout ;
wire \ShiftLeft0~54_combout ;
wire \ShiftLeft0~55_combout ;
wire \Mux26~2_combout ;
wire \ShiftRight0~52_combout ;
wire \ShiftRight0~53_combout ;
wire \ShiftRight0~54_combout ;
wire \Mux26~0_combout ;
wire \ShiftRight0~45_combout ;
wire \ShiftRight0~46_combout ;
wire \ShiftRight0~47_combout ;
wire \ShiftRight0~48_combout ;
wire \ShiftRight0~49_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftRight0~56_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~58_combout ;
wire \ShiftRight0~59_combout ;
wire \ShiftRight0~60_combout ;
wire \ShiftRight0~61_combout ;
wire \ShiftRight0~62_combout ;
wire \Mux26~1_combout ;
wire \Add0~41_combout ;
wire \Mux27~3_combout ;
wire \Mux27~4_combout ;
wire \ShiftLeft0~57_combout ;
wire \ShiftLeft0~58_combout ;
wire \ShiftLeft0~56_combout ;
wire \ShiftLeft0~59_combout ;
wire \Mux27~2_combout ;
wire \ShiftRight0~18_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~74_combout ;
wire \ShiftRight0~71_combout ;
wire \ShiftRight0~70_combout ;
wire \ShiftRight0~72_combout ;
wire \ShiftRight0~75_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftRight0~65_combout ;
wire \ShiftRight0~66_combout ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Mux6~20_combout ;
wire \Mux4~4_combout ;
wire \Add0~87_combout ;
wire \Mux4~5_combout ;
wire \ShiftRight0~76_combout ;
wire \ShiftRight0~104_combout ;
wire \ShiftLeft0~39_combout ;
wire \ShiftLeft0~40_combout ;
wire \ShiftLeft0~41_combout ;
wire \Mux4~2_combout ;
wire \ShiftLeft0~60_combout ;
wire \ShiftLeft0~61_combout ;
wire \ShiftLeft0~62_combout ;
wire \Mux4~3_combout ;
wire \Mux4~7_combout ;
wire \ShiftLeft0~64_combout ;
wire \ShiftLeft0~65_combout ;
wire \ShiftLeft0~63_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux5~7_combout ;
wire \ShiftRight0~77_combout ;
wire \ShiftRight0~105_combout ;
wire \Mux5~4_combout ;
wire \Add0~85_combout ;
wire \Mux5~5_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftLeft0~68_combout ;
wire \ShiftLeft0~69_combout ;
wire \ShiftLeft0~28_combout ;
wire \ShiftLeft0~66_combout ;
wire \ShiftLeft0~67_combout ;
wire \ShiftLeft0~70_combout ;
wire \ShiftLeft0~73_combout ;
wire \ShiftLeft0~75_combout ;
wire \Mux6~12_combout ;
wire \ShiftLeft0~76_combout ;
wire \ShiftLeft0~77_combout ;
wire \ShiftLeft0~78_combout ;
wire \ShiftLeft0~79_combout ;
wire \Mux6~13_combout ;
wire \Mux6~19_combout ;
wire \Add0~83_combout ;
wire \Mux6~14_combout ;
wire \Mux6~15_combout ;
wire \ShiftRight0~79_combout ;
wire \ShiftLeft0~85_combout ;
wire \ShiftLeft0~86_combout ;
wire \ShiftLeft0~87_combout ;
wire \ShiftLeft0~74_combout ;
wire \ShiftLeft0~84_combout ;
wire \ShiftLeft0~81_combout ;
wire \ShiftLeft0~82_combout ;
wire \ShiftLeft0~83_combout ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \Mux7~7_combout ;
wire \Mux7~4_combout ;
wire \Add0~81_combout ;
wire \Mux7~5_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Mux3~6_combout ;
wire \Mux2~0_combout ;
wire \Mux3~5_combout ;
wire \ShiftLeft0~88_combout ;
wire \Mux3~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~2_combout ;
wire \Mux3~1_combout ;
wire \ShiftLeft0~89_combout ;
wire \Mux3~2_combout ;
wire \ShiftRight0~73_combout ;
wire \ShiftRight0~80_combout ;
wire \Mux2~3_combout ;
wire \Add0~89_combout ;
wire \Mux3~3_combout ;
wire \Mux3~4_combout ;
wire \Mux2~10_combout ;
wire \ShiftLeft0~90_combout ;
wire \Mux2~5_combout ;
wire \ShiftLeft0~71_combout ;
wire \ShiftLeft0~72_combout ;
wire \ShiftLeft0~91_combout ;
wire \Mux2~7_combout ;
wire \Mux2~4_combout ;
wire \Add0~91_combout ;
wire \Mux2~8_combout ;
wire \Mux2~9_combout ;
wire \Add0~22_combout ;
wire \Add0~49_combout ;
wire \ShiftRight0~82_combout ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \Mux23~4_combout ;
wire \Mux23~5_combout ;
wire \ShiftRight0~83_combout ;
wire \Mux23~6_combout ;
wire \Add0~21_combout ;
wire \Add0~51_combout ;
wire \ShiftRight0~50_combout ;
wire \ShiftRight0~51_combout ;
wire \ShiftRight0~85_combout ;
wire \ShiftRight0~84_combout ;
wire \Mux18~4_combout ;
wire \Mux22~2_combout ;
wire \Mux22~3_combout ;
wire \Mux22~4_combout ;
wire \ShiftRight0~87_combout ;
wire \ShiftRight0~86_combout ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \Mux21~4_combout ;
wire \Add0~53_combout ;
wire \Add0~55_combout ;
wire \ShiftRight0~89_combout ;
wire \ShiftRight0~88_combout ;
wire \Mux20~2_combout ;
wire \Mux20~3_combout ;
wire \Mux20~4_combout ;
wire \Add0~18_combout ;
wire \Add0~57_combout ;
wire \Mux19~3_combout ;
wire \Mux19~4_combout ;
wire \Add0~59_combout ;
wire \ShiftRight0~81_combout ;
wire \Mux18~6_combout ;
wire \Mux18~7_combout ;
wire \Add0~61_combout ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux17~4_combout ;
wire \Add0~63_combout ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \Mux16~4_combout ;
wire \Mux29~5_combout ;
wire \Mux6~17_combout ;
wire \ShiftRight0~91_combout ;
wire \Mux28~1_combout ;
wire \Mux28~0_combout ;
wire \ShiftLeft0~92_combout ;
wire \Mux29~2_combout ;
wire \ShiftRight0~68_combout ;
wire \ShiftRight0~90_combout ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Mux29~3_combout ;
wire \Mux29~4_combout ;
wire \Mux28~6_combout ;
wire \ShiftRight0~92_combout ;
wire \ShiftRight0~19_combout ;
wire \ShiftRight0~20_combout ;
wire \Mux28~2_combout ;
wire \Mux28~3_combout ;
wire \ShiftLeft0~93_combout ;
wire \Mux28~4_combout ;
wire \ShiftRight0~93_combout ;
wire \Mux28~5_combout ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux0~7_combout ;
wire \Mux8~6_combout ;
wire \Mux8~7_combout ;
wire \Add0~79_combout ;
wire \Mux8~9_combout ;
wire \Mux15~2_combout ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \Mux10~4_combout ;
wire \Add0~9_combout ;
wire \Add0~75_combout ;
wire \Add0~8_combout ;
wire \Add0~77_combout ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux30~3_combout ;
wire \Add0~35_combout ;
wire \Mux30~4_combout ;
wire \ShiftRight0~94_combout ;
wire \ShiftRight0~95_combout ;
wire \ShiftRight0~96_combout ;
wire \ShiftRight0~97_combout ;
wire \ShiftRight0~98_combout ;
wire \ShiftRight0~99_combout ;
wire \ShiftRight0~100_combout ;
wire \Mux30~1_combout ;
wire \Mux14~8_combout ;
wire \Mux30~2_combout ;
wire \Add0~14_combout ;
wire \Add0~65_combout ;
wire \ShiftRight0~101_combout ;
wire \ShiftRight0~102_combout ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \Add0~67_combout ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \Add0~12_combout ;
wire \Add0~69_combout ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \Mux13~4_combout ;
wire \Add0~11_combout ;
wire \Add0~71_combout ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Mux12~4_combout ;
wire \Add0~10_combout ;
wire \Add0~73_combout ;
wire \Mux11~3_combout ;
wire \Mux11~4_combout ;
wire \Mux31~1_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \LessThan0~35_cout ;
wire \LessThan0~37_cout ;
wire \LessThan0~39_cout ;
wire \LessThan0~41_cout ;
wire \LessThan0~43_cout ;
wire \LessThan0~45_cout ;
wire \LessThan0~47_cout ;
wire \LessThan0~49_cout ;
wire \LessThan0~51_cout ;
wire \LessThan0~53_cout ;
wire \LessThan0~55_cout ;
wire \LessThan0~57_cout ;
wire \LessThan0~59_cout ;
wire \LessThan0~61_cout ;
wire \LessThan0~62_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~31_cout ;
wire \LessThan1~33_cout ;
wire \LessThan1~35_cout ;
wire \LessThan1~37_cout ;
wire \LessThan1~39_cout ;
wire \LessThan1~41_cout ;
wire \LessThan1~43_cout ;
wire \LessThan1~45_cout ;
wire \LessThan1~47_cout ;
wire \LessThan1~49_cout ;
wire \LessThan1~51_cout ;
wire \LessThan1~53_cout ;
wire \LessThan1~55_cout ;
wire \LessThan1~57_cout ;
wire \LessThan1~59_cout ;
wire \LessThan1~61_cout ;
wire \LessThan1~62_combout ;
wire \Mux31~2_combout ;
wire \Mux31~3_combout ;
wire \Equal0~6_combout ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \Equal0~5_combout ;
wire \Mux31~4_combout ;
wire \Mux31~5_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~69_combout ;
wire \Mux31~6_combout ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \Mux31~9_combout ;
wire \Add0~33_combout ;
wire \Mux31~10_combout ;
wire \Mux31~11_combout ;
wire \Equal0~7_combout ;
wire \Equal0~8_combout ;
wire \Equal0~9_combout ;


// Location: LCCOMB_X58_Y44_N22
cycloneive_lcell_comb \Add0~37 (
// Equation(s):
// \Add0~37_combout  = (\Add0~28_combout  & ((Mux29 & (\Add0~36  & VCC)) # (!Mux29 & (!\Add0~36 )))) # (!\Add0~28_combout  & ((Mux29 & (!\Add0~36 )) # (!Mux29 & ((\Add0~36 ) # (GND)))))
// \Add0~38  = CARRY((\Add0~28_combout  & (!Mux29 & !\Add0~36 )) # (!\Add0~28_combout  & ((!\Add0~36 ) # (!Mux29))))

	.dataa(\Add0~28_combout ),
	.datab(Mux29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~36 ),
	.combout(\Add0~37_combout ),
	.cout(\Add0~38 ));
// synopsys translate_off
defparam \Add0~37 .lut_mask = 16'h9617;
defparam \Add0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N24
cycloneive_lcell_comb \Add0~39 (
// Equation(s):
// \Add0~39_combout  = ((\Add0~27_combout  $ (Mux28 $ (!\Add0~38 )))) # (GND)
// \Add0~40  = CARRY((\Add0~27_combout  & ((Mux28) # (!\Add0~38 ))) # (!\Add0~27_combout  & (Mux28 & !\Add0~38 )))

	.dataa(\Add0~27_combout ),
	.datab(Mux28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~38 ),
	.combout(\Add0~39_combout ),
	.cout(\Add0~40 ));
// synopsys translate_off
defparam \Add0~39 .lut_mask = 16'h698E;
defparam \Add0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N4
cycloneive_lcell_comb \Add0~1 (
// Equation(s):
// \Add0~1_combout  = Selector3 $ (((\Selector71~0_combout ) # ((\Selector95~0_combout  & Mux34))))

	.dataa(Selector3),
	.datab(Selector95),
	.datac(Selector71),
	.datad(Mux34),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~1 .lut_mask = 16'h565A;
defparam \Add0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N20
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = Selector3 $ (((\Selector72~0_combout ) # ((Mux35 & \Selector95~0_combout ))))

	.dataa(Selector3),
	.datab(Mux35),
	.datac(Selector72),
	.datad(Selector95),
	.cin(gnd),
	.combout(\Add0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h565A;
defparam \Add0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N24
cycloneive_lcell_comb \Add0~3 (
// Equation(s):
// \Add0~3_combout  = Selector3 $ (((\Selector73~0_combout ) # ((Mux36 & \Selector95~0_combout ))))

	.dataa(Mux36),
	.datab(Selector73),
	.datac(Selector3),
	.datad(Selector95),
	.cin(gnd),
	.combout(\Add0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~3 .lut_mask = 16'h1E3C;
defparam \Add0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N2
cycloneive_lcell_comb \Add0~5 (
// Equation(s):
// \Add0~5_combout  = Selector3 $ (((\Selector75~0_combout ) # ((Mux38 & \Selector95~0_combout ))))

	.dataa(Selector3),
	.datab(Mux38),
	.datac(Selector95),
	.datad(Selector75),
	.cin(gnd),
	.combout(\Add0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~5 .lut_mask = 16'h556A;
defparam \Add0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N14
cycloneive_lcell_comb \Add0~7 (
// Equation(s):
// \Add0~7_combout  = Selector3 $ (((\Selector77~0_combout ) # ((Mux40 & \Selector95~0_combout ))))

	.dataa(Selector77),
	.datab(Selector3),
	.datac(Mux40),
	.datad(Selector95),
	.cin(gnd),
	.combout(\Add0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~7 .lut_mask = 16'h3666;
defparam \Add0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N14
cycloneive_lcell_comb \Add0~25 (
// Equation(s):
// \Add0~25_combout  = Selector3 $ (((\Selector95~2_combout ) # ((\Selector95~0_combout  & Mux58))))

	.dataa(Selector95),
	.datab(Selector3),
	.datac(Selector951),
	.datad(Mux58),
	.cin(gnd),
	.combout(\Add0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~25 .lut_mask = 16'h363C;
defparam \Add0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N6
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = Selector3 $ (((\Selector96~1_combout ) # ((Mux59 & \Selector100~0_combout ))))

	.dataa(Mux59),
	.datab(Selector100),
	.datac(Selector3),
	.datad(Selector96),
	.cin(gnd),
	.combout(\Add0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h0F78;
defparam \Add0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N18
cycloneive_lcell_comb \Add0~27 (
// Equation(s):
// \Add0~27_combout  = Selector3 $ (((\Selector97~1_combout ) # ((Mux60 & \Selector100~0_combout ))))

	.dataa(Mux60),
	.datab(Selector97),
	.datac(Selector100),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Add0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~27 .lut_mask = 16'h13EC;
defparam \Add0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N6
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = Selector3 $ (((\Selector98~1_combout ) # ((\Selector100~0_combout  & Mux61))))

	.dataa(Selector98),
	.datab(Selector100),
	.datac(Selector3),
	.datad(Mux61),
	.cin(gnd),
	.combout(\Add0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'h1E5A;
defparam \Add0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N12
cycloneive_lcell_comb \Add0~29 (
// Equation(s):
// \Add0~29_combout  = Selector3 $ (((\Selector99~1_combout ) # ((Mux62 & \Selector100~0_combout ))))

	.dataa(Mux62),
	.datab(Selector3),
	.datac(Selector99),
	.datad(Selector100),
	.cin(gnd),
	.combout(\Add0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~29 .lut_mask = 16'h363C;
defparam \Add0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N14
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = Selector3 $ (((\Selector100~3_combout ) # ((Mux63 & \Selector100~0_combout ))))

	.dataa(Mux63),
	.datab(Selector3),
	.datac(Selector1001),
	.datad(Selector100),
	.cin(gnd),
	.combout(\Add0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h363C;
defparam \Add0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N22
cycloneive_lcell_comb \ShiftLeft0~11 (
// Equation(s):
// \ShiftLeft0~11_combout  = (\Selector93~1_combout ) # ((\Selector92~1_combout ) # ((\Selector95~3_combout ) # (\Selector94~1_combout )))

	.dataa(Selector931),
	.datab(Selector921),
	.datac(Selector952),
	.datad(Selector941),
	.cin(gnd),
	.combout(\ShiftLeft0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~11 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N16
cycloneive_lcell_comb \ShiftRight0~37 (
// Equation(s):
// \ShiftRight0~37_combout  = (!\Selector100~4_combout  & ((\Selector99~2_combout  & (Mux23)) # (!\Selector99~2_combout  & ((Mux25)))))

	.dataa(Mux23),
	.datab(Selector991),
	.datac(Mux25),
	.datad(Selector1002),
	.cin(gnd),
	.combout(\ShiftRight0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~37 .lut_mask = 16'h00B8;
defparam \ShiftRight0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N6
cycloneive_lcell_comb \ShiftRight0~38 (
// Equation(s):
// \ShiftRight0~38_combout  = (\ShiftRight0~37_combout ) # ((\Selector100~4_combout  & \ShiftRight0~19_combout ))

	.dataa(Selector1002),
	.datab(\ShiftRight0~37_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~19_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~38 .lut_mask = 16'hEECC;
defparam \ShiftRight0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N26
cycloneive_lcell_comb \ShiftLeft0~80 (
// Equation(s):
// \ShiftLeft0~80_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~33_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~71_combout ))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftLeft0~71_combout ),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~80 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N12
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (\Mux2~2_combout  & (\ShiftLeft0~75_combout  & (!\Mux2~1_combout ))) # (!\Mux2~2_combout  & (((\Mux2~1_combout ) # (\ShiftLeft0~38_combout ))))

	.dataa(\ShiftLeft0~75_combout ),
	.datab(\Mux2~2_combout ),
	.datac(\Mux2~1_combout ),
	.datad(\ShiftLeft0~38_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'h3B38;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N22
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (\Mux0~4_combout  & ((\Selector97~2_combout  & ((\ShiftLeft0~59_combout ))) # (!\Selector97~2_combout  & (\ShiftLeft0~88_combout ))))

	.dataa(\Mux0~4_combout ),
	.datab(Selector971),
	.datac(\ShiftLeft0~88_combout ),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hA820;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N30
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (\Mux0~4_combout  & ((\Selector97~2_combout  & (\ShiftLeft0~55_combout )) # (!\Selector97~2_combout  & ((\ShiftLeft0~90_combout )))))

	.dataa(\Mux0~4_combout ),
	.datab(Selector971),
	.datac(\ShiftLeft0~55_combout ),
	.datad(\ShiftLeft0~90_combout ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hA280;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N26
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (\ShiftRight0~21_combout  & (\Mux15~2_combout  & Mux31))

	.dataa(gnd),
	.datab(\ShiftRight0~21_combout ),
	.datac(\Mux15~2_combout ),
	.datad(Mux31),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hC000;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N14
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (\ShiftLeft0~59_combout  & \Mux15~2_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~59_combout ),
	.datad(\Mux15~2_combout ),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hF000;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N30
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (\Mux15~2_combout  & ((\Selector98~2_combout  & (\ShiftLeft0~44_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~46_combout )))))

	.dataa(\ShiftLeft0~44_combout ),
	.datab(Selector981),
	.datac(\ShiftLeft0~46_combout ),
	.datad(\Mux15~2_combout ),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hB800;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N26
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (\Mux15~2_combout  & ((\Selector98~2_combout  & (\ShiftLeft0~20_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~23_combout )))))

	.dataa(\ShiftLeft0~20_combout ),
	.datab(Selector981),
	.datac(\Mux15~2_combout ),
	.datad(\ShiftLeft0~23_combout ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hB080;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N2
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// Mux110 = (\Mux23~3_combout  & ((\Add0~93_combout ) # ((\Mux23~2_combout  & \Mux1~6_combout )))) # (!\Mux23~3_combout  & (\Mux23~2_combout  & (\Mux1~6_combout )))

	.dataa(\Mux23~3_combout ),
	.datab(\Mux23~2_combout ),
	.datac(\Mux1~6_combout ),
	.datad(\Add0~93_combout ),
	.cin(gnd),
	.combout(Mux110),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hEAC0;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N22
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// Mux311 = (Selector1 & !Selector0)

	.dataa(gnd),
	.datab(Selector1),
	.datac(gnd),
	.datad(Selector0),
	.cin(gnd),
	.combout(Mux311),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'h00CC;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N12
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// Mux111 = (\Selector70~1_combout  & (Selector2 $ (((Selector3) # (Mux1))))) # (!\Selector70~1_combout  & ((Selector2 & (Selector3 $ (Mux1))) # (!Selector2 & (Selector3 & Mux1))))

	.dataa(Selector701),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Mux1),
	.cin(gnd),
	.combout(Mux111),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'h3668;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N18
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// Mux01 = (\Mux23~3_combout  & ((\Add0~96_combout ) # ((\Mux23~2_combout  & \Mux0~12_combout )))) # (!\Mux23~3_combout  & (\Mux23~2_combout  & (\Mux0~12_combout )))

	.dataa(\Mux23~3_combout ),
	.datab(\Mux23~2_combout ),
	.datac(\Mux0~12_combout ),
	.datad(\Add0~96_combout ),
	.cin(gnd),
	.combout(Mux01),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hEAC0;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N16
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// Mux02 = (Selector3 & (Selector2 $ (((Mux0) # (\Selector69~1_combout ))))) # (!Selector3 & ((Selector2 & (Mux0 $ (\Selector69~1_combout ))) # (!Selector2 & (Mux0 & \Selector69~1_combout ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(Mux0),
	.datad(Selector691),
	.cin(gnd),
	.combout(Mux02),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'h5668;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N26
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// Mux241 = (\Mux24~10_combout  & ((\Mux24~8_combout  & (\Mux24~6_combout )) # (!\Mux24~8_combout  & ((\Mux24~5_combout ))))) # (!\Mux24~10_combout  & (\Mux24~8_combout ))

	.dataa(\Mux24~10_combout ),
	.datab(\Mux24~8_combout ),
	.datac(\Mux24~6_combout ),
	.datad(\Mux24~5_combout ),
	.cin(gnd),
	.combout(Mux241),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hE6C4;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N28
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// Mux251 = (\Mux25~4_combout  & ((\Mux25~2_combout ) # ((!\Mux24~10_combout )))) # (!\Mux25~4_combout  & (((\Mux25~1_combout  & \Mux24~10_combout ))))

	.dataa(\Mux25~2_combout ),
	.datab(\Mux25~1_combout ),
	.datac(\Mux25~4_combout ),
	.datad(\Mux24~10_combout ),
	.cin(gnd),
	.combout(Mux251),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hACF0;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N18
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// Mux261 = (\Mux24~10_combout  & ((\Mux26~4_combout  & (\Mux26~2_combout )) # (!\Mux26~4_combout  & ((\Mux26~1_combout ))))) # (!\Mux24~10_combout  & (\Mux26~4_combout ))

	.dataa(\Mux24~10_combout ),
	.datab(\Mux26~4_combout ),
	.datac(\Mux26~2_combout ),
	.datad(\Mux26~1_combout ),
	.cin(gnd),
	.combout(Mux261),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hE6C4;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N24
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// Mux271 = (\Mux27~4_combout  & ((\Mux27~2_combout ) # ((!\Mux24~10_combout )))) # (!\Mux27~4_combout  & (((\Mux24~10_combout  & \Mux27~1_combout ))))

	.dataa(\Mux27~4_combout ),
	.datab(\Mux27~2_combout ),
	.datac(\Mux24~10_combout ),
	.datad(\Mux27~1_combout ),
	.cin(gnd),
	.combout(Mux271),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hDA8A;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N14
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// Mux410 = (\Mux6~20_combout  & ((\Mux4~5_combout  & ((\Mux4~7_combout ))) # (!\Mux4~5_combout  & (\ShiftRight0~104_combout )))) # (!\Mux6~20_combout  & (\Mux4~5_combout ))

	.dataa(\Mux6~20_combout ),
	.datab(\Mux4~5_combout ),
	.datac(\ShiftRight0~104_combout ),
	.datad(\Mux4~7_combout ),
	.cin(gnd),
	.combout(Mux410),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hEC64;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N30
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// Mux510 = (\Mux6~20_combout  & ((\Mux5~5_combout  & (\Mux5~7_combout )) # (!\Mux5~5_combout  & ((\ShiftRight0~105_combout ))))) # (!\Mux6~20_combout  & (((\Mux5~5_combout ))))

	.dataa(\Mux6~20_combout ),
	.datab(\Mux5~7_combout ),
	.datac(\ShiftRight0~105_combout ),
	.datad(\Mux5~5_combout ),
	.cin(gnd),
	.combout(Mux510),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hDDA0;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N0
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// Mux64 = (\Mux6~20_combout  & ((\Mux6~15_combout  & ((\Mux6~19_combout ))) # (!\Mux6~15_combout  & (\ShiftRight0~78_combout )))) # (!\Mux6~20_combout  & (((\Mux6~15_combout ))))

	.dataa(\Mux6~20_combout ),
	.datab(\ShiftRight0~78_combout ),
	.datac(\Mux6~19_combout ),
	.datad(\Mux6~15_combout ),
	.cin(gnd),
	.combout(Mux64),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hF588;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N24
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// Mux71 = (\Mux7~5_combout  & (((\Mux7~7_combout ) # (!\Mux6~20_combout )))) # (!\Mux7~5_combout  & (\ShiftRight0~79_combout  & ((\Mux6~20_combout ))))

	.dataa(\ShiftRight0~79_combout ),
	.datab(\Mux7~7_combout ),
	.datac(\Mux7~5_combout ),
	.datad(\Mux6~20_combout ),
	.cin(gnd),
	.combout(Mux71),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hCAF0;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N4
cycloneive_lcell_comb \Equal0~2 (
// Equation(s):
// Equal0 = (!Mux03 & ((Selector0) # ((!\Equal0~0_combout  & !\Equal0~1_combout ))))

	.dataa(\Equal0~0_combout ),
	.datab(Selector0),
	.datac(Mux03),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~2 .lut_mask = 16'h0C0D;
defparam \Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N12
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// Mux310 = (\Mux3~6_combout  & ((Mux311) # ((\Mux3~5_combout  & \Mux3~4_combout )))) # (!\Mux3~6_combout  & (((\Mux3~5_combout  & \Mux3~4_combout ))))

	.dataa(\Mux3~6_combout ),
	.datab(Mux311),
	.datac(\Mux3~5_combout ),
	.datad(\Mux3~4_combout ),
	.cin(gnd),
	.combout(Mux310),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hF888;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N28
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// Mux210 = (\Mux3~5_combout  & ((\Mux2~9_combout ) # ((Mux311 & \Mux2~10_combout )))) # (!\Mux3~5_combout  & (Mux311 & (\Mux2~10_combout )))

	.dataa(\Mux3~5_combout ),
	.datab(Mux311),
	.datac(\Mux2~10_combout ),
	.datad(\Mux2~9_combout ),
	.cin(gnd),
	.combout(Mux210),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hEAC0;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N22
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// Mux231 = (\Add0~49_combout  & ((\Mux23~3_combout ) # ((\Mux23~2_combout  & \Mux23~6_combout )))) # (!\Add0~49_combout  & (\Mux23~2_combout  & ((\Mux23~6_combout ))))

	.dataa(\Add0~49_combout ),
	.datab(\Mux23~2_combout ),
	.datac(\Mux23~3_combout ),
	.datad(\Mux23~6_combout ),
	.cin(gnd),
	.combout(Mux231),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hECA0;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N2
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// Mux232 = (Mux23 & (Selector2 $ (((Selector3) # (\Selector92~1_combout ))))) # (!Mux23 & ((Selector2 & (Selector3 $ (\Selector92~1_combout ))) # (!Selector2 & (Selector3 & \Selector92~1_combout ))))

	.dataa(Mux23),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector921),
	.cin(gnd),
	.combout(Mux232),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'h3668;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N18
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// Mux221 = (\Mux23~2_combout  & ((\Mux22~4_combout ) # ((\Mux23~3_combout  & \Add0~51_combout )))) # (!\Mux23~2_combout  & (\Mux23~3_combout  & (\Add0~51_combout )))

	.dataa(\Mux23~2_combout ),
	.datab(\Mux23~3_combout ),
	.datac(\Add0~51_combout ),
	.datad(\Mux22~4_combout ),
	.cin(gnd),
	.combout(Mux221),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hEAC0;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N0
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// Mux222 = (\Selector91~1_combout  & (Selector2 $ (((Selector3) # (Mux22))))) # (!\Selector91~1_combout  & ((Selector2 & (Selector3 $ (Mux22))) # (!Selector2 & (Selector3 & Mux22))))

	.dataa(Selector911),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Mux22),
	.cin(gnd),
	.combout(Mux222),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'h3668;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N22
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// Mux211 = (\Mux23~2_combout  & ((\Mux21~4_combout ) # ((\Mux23~3_combout  & \Add0~53_combout )))) # (!\Mux23~2_combout  & (\Mux23~3_combout  & ((\Add0~53_combout ))))

	.dataa(\Mux23~2_combout ),
	.datab(\Mux23~3_combout ),
	.datac(\Mux21~4_combout ),
	.datad(\Add0~53_combout ),
	.cin(gnd),
	.combout(Mux211),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hECA0;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N24
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// Mux212 = (\Selector90~1_combout  & (Selector2 $ (((Selector3) # (Mux21))))) # (!\Selector90~1_combout  & ((Selector2 & (Selector3 $ (Mux21))) # (!Selector2 & (Selector3 & Mux21))))

	.dataa(Selector901),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Mux21),
	.cin(gnd),
	.combout(Mux212),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'h3668;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N20
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// Mux201 = (\Add0~55_combout  & ((\Mux23~3_combout ) # ((\Mux23~2_combout  & \Mux20~4_combout )))) # (!\Add0~55_combout  & (\Mux23~2_combout  & ((\Mux20~4_combout ))))

	.dataa(\Add0~55_combout ),
	.datab(\Mux23~2_combout ),
	.datac(\Mux23~3_combout ),
	.datad(\Mux20~4_combout ),
	.cin(gnd),
	.combout(Mux201),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hECA0;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N10
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// Mux202 = (Mux20 & (Selector2 $ (((Selector3) # (\Selector89~1_combout ))))) # (!Mux20 & ((Selector2 & (Selector3 $ (\Selector89~1_combout ))) # (!Selector2 & (Selector3 & \Selector89~1_combout ))))

	.dataa(Mux20),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector891),
	.cin(gnd),
	.combout(Mux202),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'h3668;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N0
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// Mux191 = (\Mux23~3_combout  & ((\Add0~57_combout ) # ((\Mux23~2_combout  & \Mux19~4_combout )))) # (!\Mux23~3_combout  & (((\Mux23~2_combout  & \Mux19~4_combout ))))

	.dataa(\Mux23~3_combout ),
	.datab(\Add0~57_combout ),
	.datac(\Mux23~2_combout ),
	.datad(\Mux19~4_combout ),
	.cin(gnd),
	.combout(Mux191),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hF888;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N20
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// Mux192 = (Selector3 & (Selector2 $ (((\Selector88~1_combout ) # (Mux19))))) # (!Selector3 & ((Selector2 & (\Selector88~1_combout  $ (Mux19))) # (!Selector2 & (\Selector88~1_combout  & Mux19))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(Selector881),
	.datad(Mux19),
	.cin(gnd),
	.combout(Mux192),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'h5668;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N12
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// Mux181 = (\Mux23~3_combout  & ((\Add0~59_combout ) # ((\Mux23~2_combout  & \Mux18~7_combout )))) # (!\Mux23~3_combout  & (\Mux23~2_combout  & ((\Mux18~7_combout ))))

	.dataa(\Mux23~3_combout ),
	.datab(\Mux23~2_combout ),
	.datac(\Add0~59_combout ),
	.datad(\Mux18~7_combout ),
	.cin(gnd),
	.combout(Mux181),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hECA0;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N12
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// Mux182 = (Mux18 & (Selector2 $ (((Selector3) # (\Selector87~1_combout ))))) # (!Mux18 & ((Selector2 & (Selector3 $ (\Selector87~1_combout ))) # (!Selector2 & (Selector3 & \Selector87~1_combout ))))

	.dataa(Mux18),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector871),
	.cin(gnd),
	.combout(Mux182),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'h3668;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N28
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// Mux171 = (\Mux23~2_combout  & ((\Mux17~4_combout ) # ((\Mux23~3_combout  & \Add0~61_combout )))) # (!\Mux23~2_combout  & (\Mux23~3_combout  & (\Add0~61_combout )))

	.dataa(\Mux23~2_combout ),
	.datab(\Mux23~3_combout ),
	.datac(\Add0~61_combout ),
	.datad(\Mux17~4_combout ),
	.cin(gnd),
	.combout(Mux171),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hEAC0;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N18
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// Mux172 = (Mux17 & (Selector2 $ (((Selector3) # (\Selector86~1_combout ))))) # (!Mux17 & ((Selector2 & (Selector3 $ (\Selector86~1_combout ))) # (!Selector2 & (Selector3 & \Selector86~1_combout ))))

	.dataa(Mux17),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector861),
	.cin(gnd),
	.combout(Mux172),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'h3668;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N12
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// Mux161 = (\Mux23~3_combout  & ((\Add0~63_combout ) # ((\Mux23~2_combout  & \Mux16~4_combout )))) # (!\Mux23~3_combout  & (\Mux23~2_combout  & ((\Mux16~4_combout ))))

	.dataa(\Mux23~3_combout ),
	.datab(\Mux23~2_combout ),
	.datac(\Add0~63_combout ),
	.datad(\Mux16~4_combout ),
	.cin(gnd),
	.combout(Mux161),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hECA0;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N4
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// Mux162 = (\Selector85~1_combout  & (Selector2 $ (((Selector3) # (Mux16))))) # (!\Selector85~1_combout  & ((Selector3 & (Mux16 $ (Selector2))) # (!Selector3 & (Mux16 & Selector2))))

	.dataa(Selector851),
	.datab(Selector3),
	.datac(Mux16),
	.datad(Selector2),
	.cin(gnd),
	.combout(Mux162),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'h16E8;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N4
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// Mux291 = (Mux311 & ((\Mux29~5_combout ) # ((\Mux29~3_combout  & \Mux29~4_combout )))) # (!Mux311 & (((\Mux29~3_combout  & \Mux29~4_combout ))))

	.dataa(Mux311),
	.datab(\Mux29~5_combout ),
	.datac(\Mux29~3_combout ),
	.datad(\Mux29~4_combout ),
	.cin(gnd),
	.combout(Mux291),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hF888;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N8
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// Mux281 = (Mux311 & ((\Mux28~6_combout ) # ((\Mux29~4_combout  & \Mux28~5_combout )))) # (!Mux311 & (((\Mux29~4_combout  & \Mux28~5_combout ))))

	.dataa(Mux311),
	.datab(\Mux28~6_combout ),
	.datac(\Mux29~4_combout ),
	.datad(\Mux28~5_combout ),
	.cin(gnd),
	.combout(Mux281),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hF888;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N22
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// Mux81 = (\Mux8~5_combout ) # ((\Mux8~9_combout ) # ((\Mux23~2_combout  & \Mux8~7_combout )))

	.dataa(\Mux8~5_combout ),
	.datab(\Mux23~2_combout ),
	.datac(\Mux8~7_combout ),
	.datad(\Mux8~9_combout ),
	.cin(gnd),
	.combout(Mux81),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hFFEA;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N28
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// Mux101 = (\Mux23~3_combout  & ((\Add0~75_combout ) # ((\Mux23~2_combout  & \Mux10~4_combout )))) # (!\Mux23~3_combout  & (\Mux23~2_combout  & (\Mux10~4_combout )))

	.dataa(\Mux23~3_combout ),
	.datab(\Mux23~2_combout ),
	.datac(\Mux10~4_combout ),
	.datad(\Add0~75_combout ),
	.cin(gnd),
	.combout(Mux101),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hEAC0;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N28
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// Mux102 = (\Selector79~1_combout  & (Selector2 $ (((Mux10) # (Selector3))))) # (!\Selector79~1_combout  & ((Mux10 & (Selector3 $ (Selector2))) # (!Mux10 & (Selector3 & Selector2))))

	.dataa(Selector791),
	.datab(Mux10),
	.datac(Selector3),
	.datad(Selector2),
	.cin(gnd),
	.combout(Mux102),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'h16E8;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N18
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// Mux91 = (\Mux23~3_combout  & ((\Add0~77_combout ) # ((\Mux23~2_combout  & \Mux9~5_combout )))) # (!\Mux23~3_combout  & (((\Mux23~2_combout  & \Mux9~5_combout ))))

	.dataa(\Mux23~3_combout ),
	.datab(\Add0~77_combout ),
	.datac(\Mux23~2_combout ),
	.datad(\Mux9~5_combout ),
	.cin(gnd),
	.combout(Mux91),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hF888;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N6
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// Mux92 = (Mux9 & (Selector2 $ (((Selector3) # (\Selector78~1_combout ))))) # (!Mux9 & ((Selector2 & (Selector3 $ (\Selector78~1_combout ))) # (!Selector2 & (Selector3 & \Selector78~1_combout ))))

	.dataa(Mux9),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector781),
	.cin(gnd),
	.combout(Mux92),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'h3668;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N6
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// Mux301 = (!Selector0 & ((\Mux30~4_combout ) # ((\Mux30~1_combout ) # (\Mux30~2_combout ))))

	.dataa(Selector0),
	.datab(\Mux30~4_combout ),
	.datac(\Mux30~1_combout ),
	.datad(\Mux30~2_combout ),
	.cin(gnd),
	.combout(Mux301),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'h5554;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N0
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// Mux151 = (\Mux23~2_combout  & ((\Mux15~5_combout ) # ((\Mux23~3_combout  & \Add0~65_combout )))) # (!\Mux23~2_combout  & (\Mux23~3_combout  & (\Add0~65_combout )))

	.dataa(\Mux23~2_combout ),
	.datab(\Mux23~3_combout ),
	.datac(\Add0~65_combout ),
	.datad(\Mux15~5_combout ),
	.cin(gnd),
	.combout(Mux151),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hEAC0;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N28
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// Mux152 = (Mux15 & (Selector2 $ (((Selector3) # (\Selector84~2_combout ))))) # (!Mux15 & ((Selector2 & (Selector3 $ (\Selector84~2_combout ))) # (!Selector2 & (Selector3 & \Selector84~2_combout ))))

	.dataa(Mux15),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector841),
	.cin(gnd),
	.combout(Mux152),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'h3668;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N8
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// Mux141 = (\Mux23~2_combout  & ((\Mux14~5_combout ) # ((\Mux23~3_combout  & \Add0~67_combout )))) # (!\Mux23~2_combout  & (\Mux23~3_combout  & (\Add0~67_combout )))

	.dataa(\Mux23~2_combout ),
	.datab(\Mux23~3_combout ),
	.datac(\Add0~67_combout ),
	.datad(\Mux14~5_combout ),
	.cin(gnd),
	.combout(Mux141),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hEAC0;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N26
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// Mux142 = (\Selector83~1_combout  & (Selector2 $ (((Selector3) # (Mux14))))) # (!\Selector83~1_combout  & ((Selector3 & (Mux14 $ (Selector2))) # (!Selector3 & (Mux14 & Selector2))))

	.dataa(Selector831),
	.datab(Selector3),
	.datac(Mux14),
	.datad(Selector2),
	.cin(gnd),
	.combout(Mux142),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'h16E8;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N12
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// Mux131 = (\Mux23~2_combout  & ((\Mux13~4_combout ) # ((\Mux23~3_combout  & \Add0~69_combout )))) # (!\Mux23~2_combout  & (\Mux23~3_combout  & (\Add0~69_combout )))

	.dataa(\Mux23~2_combout ),
	.datab(\Mux23~3_combout ),
	.datac(\Add0~69_combout ),
	.datad(\Mux13~4_combout ),
	.cin(gnd),
	.combout(Mux131),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hEAC0;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N10
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// Mux132 = (Selector3 & (Selector2 $ (((Mux13) # (\Selector82~1_combout ))))) # (!Selector3 & ((Selector2 & (Mux13 $ (\Selector82~1_combout ))) # (!Selector2 & (Mux13 & \Selector82~1_combout ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(Mux13),
	.datad(Selector821),
	.cin(gnd),
	.combout(Mux132),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'h5668;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N22
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// Mux121 = (\Mux23~3_combout  & ((\Add0~71_combout ) # ((\Mux23~2_combout  & \Mux12~4_combout )))) # (!\Mux23~3_combout  & (((\Mux23~2_combout  & \Mux12~4_combout ))))

	.dataa(\Mux23~3_combout ),
	.datab(\Add0~71_combout ),
	.datac(\Mux23~2_combout ),
	.datad(\Mux12~4_combout ),
	.cin(gnd),
	.combout(Mux121),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hF888;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N18
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// Mux122 = (\Selector81~1_combout  & (Selector2 $ (((Selector3) # (Mux12))))) # (!\Selector81~1_combout  & ((Selector2 & (Selector3 $ (Mux12))) # (!Selector2 & (Selector3 & Mux12))))

	.dataa(Selector811),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Mux12),
	.cin(gnd),
	.combout(Mux122),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'h3668;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N0
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// Mux112 = (\Mux23~2_combout  & ((\Mux11~4_combout ) # ((\Mux23~3_combout  & \Add0~73_combout )))) # (!\Mux23~2_combout  & (\Mux23~3_combout  & (\Add0~73_combout )))

	.dataa(\Mux23~2_combout ),
	.datab(\Mux23~3_combout ),
	.datac(\Add0~73_combout ),
	.datad(\Mux11~4_combout ),
	.cin(gnd),
	.combout(Mux112),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hEAC0;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N8
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// Mux113 = (Mux11 & (Selector2 $ (((Selector3) # (\Selector80~1_combout ))))) # (!Mux11 & ((Selector3 & (Selector2 $ (\Selector80~1_combout ))) # (!Selector3 & (Selector2 & \Selector80~1_combout ))))

	.dataa(Mux11),
	.datab(Selector3),
	.datac(Selector2),
	.datad(Selector801),
	.cin(gnd),
	.combout(Mux113),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'h1E68;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N18
cycloneive_lcell_comb \Equal0~10 (
// Equation(s):
// Equal01 = (!\Mux31~2_combout  & (!Mux210 & (!Mux310 & \Equal0~9_combout )))

	.dataa(\Mux31~2_combout ),
	.datab(Mux210),
	.datac(Mux310),
	.datad(\Equal0~9_combout ),
	.cin(gnd),
	.combout(Equal01),
	.cout());
// synopsys translate_off
defparam \Equal0~10 .lut_mask = 16'h0100;
defparam \Equal0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N26
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// Mux312 = (\Mux31~11_combout ) # ((\Mux31~2_combout ) # ((Mux311 & \Mux31~3_combout )))

	.dataa(Mux311),
	.datab(\Mux31~3_combout ),
	.datac(\Mux31~11_combout ),
	.datad(\Mux31~2_combout ),
	.cin(gnd),
	.combout(Mux312),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hFFF8;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N2
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// Mux114 = (Mux110) # ((Mux111 & (!Selector0 & Selector1)))

	.dataa(Mux111),
	.datab(Selector0),
	.datac(Selector1),
	.datad(Mux110),
	.cin(gnd),
	.combout(Mux114),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hFF20;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N10
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// Mux03 = (Mux01) # ((Selector1 & (Mux02 & !Selector0)))

	.dataa(Selector1),
	.datab(Mux02),
	.datac(Selector0),
	.datad(Mux01),
	.cin(gnd),
	.combout(Mux03),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hFF08;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N14
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// Mux233 = (Mux231) # ((Selector1 & (Mux232 & !Selector0)))

	.dataa(Selector1),
	.datab(Mux232),
	.datac(Mux231),
	.datad(Selector0),
	.cin(gnd),
	.combout(Mux233),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hF0F8;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N14
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// Mux223 = (Mux221) # ((Selector1 & (Mux222 & !Selector0)))

	.dataa(Selector1),
	.datab(Mux222),
	.datac(Selector0),
	.datad(Mux221),
	.cin(gnd),
	.combout(Mux223),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hFF08;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N16
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// Mux213 = (Mux211) # ((Selector1 & (!Selector0 & Mux212)))

	.dataa(Selector1),
	.datab(Selector0),
	.datac(Mux211),
	.datad(Mux212),
	.cin(gnd),
	.combout(Mux213),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hF2F0;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N0
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// Mux203 = (Mux201) # ((!Selector0 & (Mux202 & Selector1)))

	.dataa(Selector0),
	.datab(Mux202),
	.datac(Selector1),
	.datad(Mux201),
	.cin(gnd),
	.combout(Mux203),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hFF40;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N26
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// Mux193 = (Mux191) # ((!Selector0 & (Selector1 & Mux192)))

	.dataa(Selector0),
	.datab(Selector1),
	.datac(Mux192),
	.datad(Mux191),
	.cin(gnd),
	.combout(Mux193),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hFF40;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N22
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// Mux183 = (Mux181) # ((Mux182 & (!Selector0 & Selector1)))

	.dataa(Mux182),
	.datab(Selector0),
	.datac(Selector1),
	.datad(Mux181),
	.cin(gnd),
	.combout(Mux183),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hFF20;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N26
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// Mux173 = (Mux171) # ((!Selector0 & (Mux172 & Selector1)))

	.dataa(Selector0),
	.datab(Mux172),
	.datac(Selector1),
	.datad(Mux171),
	.cin(gnd),
	.combout(Mux173),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hFF40;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N26
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// Mux163 = (Mux161) # ((!Selector0 & (Mux162 & Selector1)))

	.dataa(Selector0),
	.datab(Mux162),
	.datac(Selector1),
	.datad(Mux161),
	.cin(gnd),
	.combout(Mux163),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hFF40;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N0
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// Mux103 = (Mux101) # ((Selector1 & (Mux102 & !Selector0)))

	.dataa(Selector1),
	.datab(Mux102),
	.datac(Selector0),
	.datad(Mux101),
	.cin(gnd),
	.combout(Mux103),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hFF08;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N6
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// Mux93 = (Mux91) # ((Mux92 & (!Selector0 & Selector1)))

	.dataa(Mux92),
	.datab(Selector0),
	.datac(Selector1),
	.datad(Mux91),
	.cin(gnd),
	.combout(Mux93),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hFF20;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N16
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// Mux153 = (Mux151) # ((Selector1 & (!Selector0 & Mux152)))

	.dataa(Selector1),
	.datab(Selector0),
	.datac(Mux152),
	.datad(Mux151),
	.cin(gnd),
	.combout(Mux153),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hFF20;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N14
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// Mux143 = (Mux141) # ((Selector1 & (!Selector0 & Mux142)))

	.dataa(Selector1),
	.datab(Selector0),
	.datac(Mux141),
	.datad(Mux142),
	.cin(gnd),
	.combout(Mux143),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hF2F0;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N24
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// Mux133 = (Mux131) # ((Selector1 & (!Selector0 & Mux132)))

	.dataa(Selector1),
	.datab(Selector0),
	.datac(Mux132),
	.datad(Mux131),
	.cin(gnd),
	.combout(Mux133),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hFF20;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N22
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// Mux123 = (Mux121) # ((Selector1 & (!Selector0 & Mux122)))

	.dataa(Selector1),
	.datab(Selector0),
	.datac(Mux122),
	.datad(Mux121),
	.cin(gnd),
	.combout(Mux123),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hFF20;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N28
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// Mux115 = (Mux112) # ((Selector1 & (!Selector0 & Mux113)))

	.dataa(Selector1),
	.datab(Selector0),
	.datac(Mux113),
	.datad(Mux112),
	.cin(gnd),
	.combout(Mux115),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hFF20;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N6
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (!Selector0 & (!Selector1 & Selector2))

	.dataa(Selector0),
	.datab(gnd),
	.datac(Selector1),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'h0500;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N24
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (!Selector2 & (!Selector1 & !Selector0))

	.dataa(Selector2),
	.datab(Selector1),
	.datac(gnd),
	.datad(Selector0),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'h0011;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N0
cycloneive_lcell_comb \ShiftLeft0~17 (
// Equation(s):
// \ShiftLeft0~17_combout  = (\Selector72~1_combout ) # ((\Selector74~1_combout ) # ((\Selector73~1_combout ) # (\Selector75~1_combout )))

	.dataa(Selector721),
	.datab(Selector741),
	.datac(Selector731),
	.datad(Selector751),
	.cin(gnd),
	.combout(\ShiftLeft0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~17 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N22
cycloneive_lcell_comb \ShiftLeft0~18 (
// Equation(s):
// \ShiftLeft0~18_combout  = (\Selector69~1_combout ) # ((\Selector71~1_combout ) # ((\Selector70~1_combout ) # (\ShiftLeft0~17_combout )))

	.dataa(Selector691),
	.datab(Selector711),
	.datac(Selector701),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~18 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N2
cycloneive_lcell_comb \ShiftLeft0~16 (
// Equation(s):
// \ShiftLeft0~16_combout  = (\Selector76~1_combout ) # ((\Selector78~1_combout ) # ((\Selector77~1_combout ) # (\Selector79~1_combout )))

	.dataa(Selector761),
	.datab(Selector781),
	.datac(Selector771),
	.datad(Selector791),
	.cin(gnd),
	.combout(\ShiftLeft0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~16 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N26
cycloneive_lcell_comb \ShiftLeft0~12 (
// Equation(s):
// \ShiftLeft0~12_combout  = (\Selector90~1_combout ) # ((\Selector89~1_combout ) # ((\Selector88~1_combout ) # (\Selector91~1_combout )))

	.dataa(Selector901),
	.datab(Selector891),
	.datac(Selector881),
	.datad(Selector911),
	.cin(gnd),
	.combout(\ShiftLeft0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~12 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N22
cycloneive_lcell_comb \ShiftLeft0~14 (
// Equation(s):
// \ShiftLeft0~14_combout  = (\Selector81~1_combout ) # ((\Selector82~1_combout ) # ((\Selector80~1_combout ) # (\Selector83~1_combout )))

	.dataa(Selector811),
	.datab(Selector821),
	.datac(Selector801),
	.datad(Selector831),
	.cin(gnd),
	.combout(\ShiftLeft0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~14 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N28
cycloneive_lcell_comb \ShiftLeft0~13 (
// Equation(s):
// \ShiftLeft0~13_combout  = (\Selector87~1_combout ) # ((\Selector86~1_combout ) # ((\Selector85~1_combout ) # (\Selector84~2_combout )))

	.dataa(Selector871),
	.datab(Selector861),
	.datac(Selector851),
	.datad(Selector841),
	.cin(gnd),
	.combout(\ShiftLeft0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~13 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N12
cycloneive_lcell_comb \ShiftLeft0~15 (
// Equation(s):
// \ShiftLeft0~15_combout  = (\ShiftLeft0~11_combout ) # ((\ShiftLeft0~12_combout ) # ((\ShiftLeft0~14_combout ) # (\ShiftLeft0~13_combout )))

	.dataa(\ShiftLeft0~11_combout ),
	.datab(\ShiftLeft0~12_combout ),
	.datac(\ShiftLeft0~14_combout ),
	.datad(\ShiftLeft0~13_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~15 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N30
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (!\Selector96~2_combout  & (!\ShiftLeft0~18_combout  & (!\ShiftLeft0~16_combout  & !\ShiftLeft0~15_combout )))

	.dataa(Selector961),
	.datab(\ShiftLeft0~18_combout ),
	.datac(\ShiftLeft0~16_combout ),
	.datad(\ShiftLeft0~15_combout ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'h0001;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N26
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (Selector3) # (!\Mux0~4_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector3),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hF0FF;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N20
cycloneive_lcell_comb \ShiftLeft0~4 (
// Equation(s):
// \ShiftLeft0~4_combout  = (\Selector99~2_combout  & (Mux11)) # (!\Selector99~2_combout  & ((Mux9)))

	.dataa(Selector991),
	.datab(gnd),
	.datac(Mux11),
	.datad(Mux9),
	.cin(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~4 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N2
cycloneive_lcell_comb \ShiftLeft0~3 (
// Equation(s):
// \ShiftLeft0~3_combout  = (\Selector99~2_combout  & ((Mux12))) # (!\Selector99~2_combout  & (Mux10))

	.dataa(Selector991),
	.datab(gnd),
	.datac(Mux10),
	.datad(Mux12),
	.cin(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~3 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N14
cycloneive_lcell_comb \ShiftLeft0~5 (
// Equation(s):
// \ShiftLeft0~5_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~3_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~4_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~4_combout ),
	.datac(Selector1002),
	.datad(\ShiftLeft0~3_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~5 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N20
cycloneive_lcell_comb \ShiftLeft0~1 (
// Equation(s):
// \ShiftLeft0~1_combout  = (\Selector99~2_combout  & ((Mux15))) # (!\Selector99~2_combout  & (Mux13))

	.dataa(Selector991),
	.datab(gnd),
	.datac(Mux13),
	.datad(Mux15),
	.cin(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~1 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N28
cycloneive_lcell_comb \ShiftLeft0~0 (
// Equation(s):
// \ShiftLeft0~0_combout  = (\Selector99~2_combout  & ((Mux16))) # (!\Selector99~2_combout  & (Mux14))

	.dataa(Selector991),
	.datab(Mux14),
	.datac(Mux16),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~0 .lut_mask = 16'hE4E4;
defparam \ShiftLeft0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N10
cycloneive_lcell_comb \ShiftLeft0~2 (
// Equation(s):
// \ShiftLeft0~2_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~0_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~1_combout ))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftLeft0~1_combout ),
	.datad(\ShiftLeft0~0_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~2 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N12
cycloneive_lcell_comb \ShiftLeft0~6 (
// Equation(s):
// \ShiftLeft0~6_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~2_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~5_combout ))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~5_combout ),
	.datad(\ShiftLeft0~2_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~6 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N0
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (\Selector98~2_combout ) # ((!\Selector99~2_combout  & \Selector100~4_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(Selector991),
	.datad(Selector1002),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hCFCC;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N22
cycloneive_lcell_comb \ShiftLeft0~8 (
// Equation(s):
// \ShiftLeft0~8_combout  = (\Selector99~2_combout  & ((\Selector100~4_combout  & ((Mux8))) # (!\Selector100~4_combout  & (Mux7))))

	.dataa(Selector1002),
	.datab(Selector991),
	.datac(Mux7),
	.datad(Mux8),
	.cin(gnd),
	.combout(\ShiftLeft0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~8 .lut_mask = 16'hC840;
defparam \ShiftLeft0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N24
cycloneive_lcell_comb \ShiftLeft0~9 (
// Equation(s):
// \ShiftLeft0~9_combout  = (\Selector100~4_combout  & ((Mux6))) # (!\Selector100~4_combout  & (Mux5))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(Mux5),
	.datad(Mux6),
	.cin(gnd),
	.combout(\ShiftLeft0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~9 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N26
cycloneive_lcell_comb \ShiftLeft0~10 (
// Equation(s):
// \ShiftLeft0~10_combout  = (\ShiftLeft0~8_combout ) # ((!\Selector99~2_combout  & \ShiftLeft0~9_combout ))

	.dataa(Selector991),
	.datab(gnd),
	.datac(\ShiftLeft0~8_combout ),
	.datad(\ShiftLeft0~9_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~10 .lut_mask = 16'hF5F0;
defparam \ShiftLeft0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N30
cycloneive_lcell_comb \ShiftLeft0~7 (
// Equation(s):
// \ShiftLeft0~7_combout  = (\Selector100~4_combout  & (Mux4)) # (!\Selector100~4_combout  & ((Mux3)))

	.dataa(Mux4),
	.datab(Selector1002),
	.datac(gnd),
	.datad(Mux3),
	.cin(gnd),
	.combout(\ShiftLeft0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~7 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N0
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (\Mux0~3_combout  & (Mux1 & ((!\Mux0~2_combout )))) # (!\Mux0~3_combout  & (((\ShiftLeft0~7_combout ) # (\Mux0~2_combout ))))

	.dataa(\Mux0~3_combout ),
	.datab(Mux1),
	.datac(\ShiftLeft0~7_combout ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'h55D8;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N16
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (\Mux0~2_combout  & ((\Mux1~2_combout  & ((\ShiftLeft0~10_combout ))) # (!\Mux1~2_combout  & (Mux2)))) # (!\Mux0~2_combout  & (((\Mux1~2_combout ))))

	.dataa(Mux2),
	.datab(\Mux0~2_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\Mux1~2_combout ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hF388;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N10
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = Selector3 $ (!\Mux0~4_combout )

	.dataa(gnd),
	.datab(Selector3),
	.datac(\Mux0~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hC3C3;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N18
cycloneive_lcell_comb \ShiftLeft0~22 (
// Equation(s):
// \ShiftLeft0~22_combout  = (\Selector99~2_combout  & (Mux27)) # (!\Selector99~2_combout  & ((Mux25)))

	.dataa(gnd),
	.datab(Selector991),
	.datac(Mux27),
	.datad(Mux25),
	.cin(gnd),
	.combout(\ShiftLeft0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~22 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N16
cycloneive_lcell_comb \ShiftLeft0~23 (
// Equation(s):
// \ShiftLeft0~23_combout  = (\Selector100~4_combout  & (\ShiftLeft0~21_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~22_combout )))

	.dataa(\ShiftLeft0~21_combout ),
	.datab(gnd),
	.datac(Selector1002),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~23 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N4
cycloneive_lcell_comb \ShiftLeft0~19 (
// Equation(s):
// \ShiftLeft0~19_combout  = (!\Selector100~4_combout  & ((\Selector99~2_combout  & ((Mux31))) # (!\Selector99~2_combout  & (Mux29))))

	.dataa(Mux29),
	.datab(Mux31),
	.datac(Selector1002),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftLeft0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~19 .lut_mask = 16'h0C0A;
defparam \ShiftLeft0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N30
cycloneive_lcell_comb \ShiftLeft0~20 (
// Equation(s):
// \ShiftLeft0~20_combout  = (\ShiftLeft0~19_combout ) # ((\Selector100~4_combout  & (Mux30 & !\Selector99~2_combout )))

	.dataa(Selector1002),
	.datab(Mux30),
	.datac(Selector991),
	.datad(\ShiftLeft0~19_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~20 .lut_mask = 16'hFF08;
defparam \ShiftLeft0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N16
cycloneive_lcell_comb \ShiftLeft0~24 (
// Equation(s):
// \ShiftLeft0~24_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~20_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~23_combout ))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~23_combout ),
	.datad(\ShiftLeft0~20_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~24 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N24
cycloneive_lcell_comb \ShiftLeft0~29 (
// Equation(s):
// \ShiftLeft0~29_combout  = (\Selector99~2_combout  & (Mux19)) # (!\Selector99~2_combout  & ((Mux17)))

	.dataa(Selector991),
	.datab(gnd),
	.datac(Mux19),
	.datad(Mux17),
	.cin(gnd),
	.combout(\ShiftLeft0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~29 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N2
cycloneive_lcell_comb \ShiftLeft0~30 (
// Equation(s):
// \ShiftLeft0~30_combout  = (\Selector100~4_combout  & (\ShiftLeft0~28_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~29_combout )))

	.dataa(\ShiftLeft0~28_combout ),
	.datab(gnd),
	.datac(Selector1002),
	.datad(\ShiftLeft0~29_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~30 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N14
cycloneive_lcell_comb \ShiftLeft0~25 (
// Equation(s):
// \ShiftLeft0~25_combout  = (\Selector99~2_combout  & (Mux24)) # (!\Selector99~2_combout  & ((Mux22)))

	.dataa(Selector991),
	.datab(gnd),
	.datac(Mux24),
	.datad(Mux22),
	.cin(gnd),
	.combout(\ShiftLeft0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~25 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N26
cycloneive_lcell_comb \ShiftLeft0~26 (
// Equation(s):
// \ShiftLeft0~26_combout  = (\Selector99~2_combout  & (Mux23)) # (!\Selector99~2_combout  & ((Mux21)))

	.dataa(Mux23),
	.datab(gnd),
	.datac(Mux21),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftLeft0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~26 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N20
cycloneive_lcell_comb \ShiftLeft0~27 (
// Equation(s):
// \ShiftLeft0~27_combout  = (\Selector100~4_combout  & (\ShiftLeft0~25_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~26_combout )))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftLeft0~25_combout ),
	.datad(\ShiftLeft0~26_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~27 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N22
cycloneive_lcell_comb \ShiftLeft0~31 (
// Equation(s):
// \ShiftLeft0~31_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~27_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~30_combout ))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~30_combout ),
	.datad(\ShiftLeft0~27_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~31 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N24
cycloneive_lcell_comb \ShiftLeft0~32 (
// Equation(s):
// \ShiftLeft0~32_combout  = (\ShiftLeft0~18_combout ) # ((\ShiftLeft0~16_combout ) # (\ShiftLeft0~15_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~18_combout ),
	.datac(\ShiftLeft0~16_combout ),
	.datad(\ShiftLeft0~15_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~32 .lut_mask = 16'hFFFC;
defparam \ShiftLeft0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N8
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (!\ShiftLeft0~32_combout  & ((\Selector97~2_combout  & (\ShiftLeft0~24_combout )) # (!\Selector97~2_combout  & ((\ShiftLeft0~31_combout )))))

	.dataa(Selector971),
	.datab(\ShiftLeft0~24_combout ),
	.datac(\ShiftLeft0~31_combout ),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'h00D8;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N0
cycloneive_lcell_comb \ShiftRight0~6 (
// Equation(s):
// \ShiftRight0~6_combout  = (\Selector100~4_combout  & ((Mux0))) # (!\Selector100~4_combout  & (Mux1))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(Mux1),
	.datad(Mux0),
	.cin(gnd),
	.combout(\ShiftRight0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~6 .lut_mask = 16'hFC30;
defparam \ShiftRight0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N22
cycloneive_lcell_comb \ShiftRight0~103 (
// Equation(s):
// \ShiftRight0~103_combout  = (!\Selector99~2_combout  & (!\Selector98~2_combout  & (\ShiftRight0~6_combout  & !\Selector97~2_combout )))

	.dataa(Selector991),
	.datab(Selector981),
	.datac(\ShiftRight0~6_combout ),
	.datad(Selector971),
	.cin(gnd),
	.combout(\ShiftRight0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~103 .lut_mask = 16'h0010;
defparam \ShiftRight0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N10
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (\Mux0~7_combout  & (\Mux0~6_combout  & ((\ShiftRight0~103_combout )))) # (!\Mux0~7_combout  & (((\Mux1~4_combout )) # (!\Mux0~6_combout )))

	.dataa(\Mux0~7_combout ),
	.datab(\Mux0~6_combout ),
	.datac(\Mux1~4_combout ),
	.datad(\ShiftRight0~103_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hD951;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N4
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (\Mux0~5_combout  & (((\Mux1~5_combout )))) # (!\Mux0~5_combout  & ((\Mux1~5_combout  & ((\Mux1~3_combout ))) # (!\Mux1~5_combout  & (\ShiftLeft0~6_combout ))))

	.dataa(\Mux0~5_combout ),
	.datab(\ShiftLeft0~6_combout ),
	.datac(\Mux1~3_combout ),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hFA44;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N30
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = Selector3 $ (((\Selector70~0_combout ) # ((\Selector95~0_combout  & Mux33))))

	.dataa(Selector70),
	.datab(Selector3),
	.datac(Selector95),
	.datad(Mux33),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h3666;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N20
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = Selector3 $ (((\Selector74~0_combout ) # ((\Selector95~0_combout  & Mux37))))

	.dataa(Selector95),
	.datab(Mux37),
	.datac(Selector3),
	.datad(Selector74),
	.cin(gnd),
	.combout(\Add0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h0F78;
defparam \Add0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N24
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = Selector3 $ (((\Selector76~0_combout ) # ((\Selector95~0_combout  & Mux39))))

	.dataa(Selector95),
	.datab(Mux39),
	.datac(Selector3),
	.datad(Selector76),
	.cin(gnd),
	.combout(\Add0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h0F78;
defparam \Add0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N10
cycloneive_lcell_comb \Add0~13 (
// Equation(s):
// \Add0~13_combout  = Selector3 $ (((\Selector83~0_combout ) # ((\Selector95~0_combout  & Mux46))))

	.dataa(Selector3),
	.datab(Selector83),
	.datac(Selector95),
	.datad(Mux46),
	.cin(gnd),
	.combout(\Add0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~13 .lut_mask = 16'h5666;
defparam \Add0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N0
cycloneive_lcell_comb \Add0~15 (
// Equation(s):
// \Add0~15_combout  = Selector3 $ (((\Selector85~0_combout ) # ((\Selector95~0_combout  & Mux48))))

	.dataa(Selector85),
	.datab(Selector95),
	.datac(Selector3),
	.datad(Mux48),
	.cin(gnd),
	.combout(\Add0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~15 .lut_mask = 16'h1E5A;
defparam \Add0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N8
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = Selector3 $ (((\Selector86~0_combout ) # ((\Selector95~0_combout  & Mux49))))

	.dataa(Selector95),
	.datab(Mux49),
	.datac(Selector3),
	.datad(Selector86),
	.cin(gnd),
	.combout(\Add0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h0F78;
defparam \Add0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N14
cycloneive_lcell_comb \Add0~17 (
// Equation(s):
// \Add0~17_combout  = Selector3 $ (((\Selector87~0_combout ) # ((Mux50 & \Selector95~0_combout ))))

	.dataa(Selector3),
	.datab(Mux50),
	.datac(Selector87),
	.datad(Selector95),
	.cin(gnd),
	.combout(\Add0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~17 .lut_mask = 16'h565A;
defparam \Add0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N30
cycloneive_lcell_comb \Add0~19 (
// Equation(s):
// \Add0~19_combout  = Selector3 $ (((\Selector89~0_combout ) # ((Mux52 & \Selector95~0_combout ))))

	.dataa(Selector3),
	.datab(Mux52),
	.datac(Selector95),
	.datad(Selector89),
	.cin(gnd),
	.combout(\Add0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~19 .lut_mask = 16'h556A;
defparam \Add0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N28
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = Selector3 $ (((\Selector90~0_combout ) # ((\Selector95~0_combout  & Mux53))))

	.dataa(Selector95),
	.datab(Mux53),
	.datac(Selector3),
	.datad(Selector90),
	.cin(gnd),
	.combout(\Add0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h0F78;
defparam \Add0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N12
cycloneive_lcell_comb \Add0~23 (
// Equation(s):
// \Add0~23_combout  = Selector3 $ (((\Selector93~0_combout ) # ((\Selector95~0_combout  & Mux56))))

	.dataa(Selector3),
	.datab(Selector95),
	.datac(Mux56),
	.datad(Selector93),
	.cin(gnd),
	.combout(\Add0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~23 .lut_mask = 16'h556A;
defparam \Add0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N4
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = Selector3 $ (((\Selector94~0_combout ) # ((\Selector95~0_combout  & Mux57))))

	.dataa(Selector95),
	.datab(Selector3),
	.datac(Mux57),
	.datad(Selector94),
	.cin(gnd),
	.combout(\Add0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'h336C;
defparam \Add0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N16
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_cout  = CARRY(Selector3)

	.dataa(gnd),
	.datab(Selector3),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add0~32_cout ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'h00CC;
defparam \Add0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N18
cycloneive_lcell_comb \Add0~33 (
// Equation(s):
// \Add0~33_combout  = (\Add0~30_combout  & ((Mux31 & (\Add0~32_cout  & VCC)) # (!Mux31 & (!\Add0~32_cout )))) # (!\Add0~30_combout  & ((Mux31 & (!\Add0~32_cout )) # (!Mux31 & ((\Add0~32_cout ) # (GND)))))
// \Add0~34  = CARRY((\Add0~30_combout  & (!Mux31 & !\Add0~32_cout )) # (!\Add0~30_combout  & ((!\Add0~32_cout ) # (!Mux31))))

	.dataa(\Add0~30_combout ),
	.datab(Mux31),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~32_cout ),
	.combout(\Add0~33_combout ),
	.cout(\Add0~34 ));
// synopsys translate_off
defparam \Add0~33 .lut_mask = 16'h9617;
defparam \Add0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N20
cycloneive_lcell_comb \Add0~35 (
// Equation(s):
// \Add0~35_combout  = ((\Add0~29_combout  $ (Mux30 $ (!\Add0~34 )))) # (GND)
// \Add0~36  = CARRY((\Add0~29_combout  & ((Mux30) # (!\Add0~34 ))) # (!\Add0~29_combout  & (Mux30 & !\Add0~34 )))

	.dataa(\Add0~29_combout ),
	.datab(Mux30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~34 ),
	.combout(\Add0~35_combout ),
	.cout(\Add0~36 ));
// synopsys translate_off
defparam \Add0~35 .lut_mask = 16'h698E;
defparam \Add0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N26
cycloneive_lcell_comb \Add0~41 (
// Equation(s):
// \Add0~41_combout  = (\Add0~26_combout  & ((Mux27 & (\Add0~40  & VCC)) # (!Mux27 & (!\Add0~40 )))) # (!\Add0~26_combout  & ((Mux27 & (!\Add0~40 )) # (!Mux27 & ((\Add0~40 ) # (GND)))))
// \Add0~42  = CARRY((\Add0~26_combout  & (!Mux27 & !\Add0~40 )) # (!\Add0~26_combout  & ((!\Add0~40 ) # (!Mux27))))

	.dataa(\Add0~26_combout ),
	.datab(Mux27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~40 ),
	.combout(\Add0~41_combout ),
	.cout(\Add0~42 ));
// synopsys translate_off
defparam \Add0~41 .lut_mask = 16'h9617;
defparam \Add0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N28
cycloneive_lcell_comb \Add0~43 (
// Equation(s):
// \Add0~43_combout  = ((\Add0~25_combout  $ (Mux26 $ (!\Add0~42 )))) # (GND)
// \Add0~44  = CARRY((\Add0~25_combout  & ((Mux26) # (!\Add0~42 ))) # (!\Add0~25_combout  & (Mux26 & !\Add0~42 )))

	.dataa(\Add0~25_combout ),
	.datab(Mux26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~42 ),
	.combout(\Add0~43_combout ),
	.cout(\Add0~44 ));
// synopsys translate_off
defparam \Add0~43 .lut_mask = 16'h698E;
defparam \Add0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N30
cycloneive_lcell_comb \Add0~45 (
// Equation(s):
// \Add0~45_combout  = (Mux25 & ((\Add0~24_combout  & (\Add0~44  & VCC)) # (!\Add0~24_combout  & (!\Add0~44 )))) # (!Mux25 & ((\Add0~24_combout  & (!\Add0~44 )) # (!\Add0~24_combout  & ((\Add0~44 ) # (GND)))))
// \Add0~46  = CARRY((Mux25 & (!\Add0~24_combout  & !\Add0~44 )) # (!Mux25 & ((!\Add0~44 ) # (!\Add0~24_combout ))))

	.dataa(Mux25),
	.datab(\Add0~24_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~44 ),
	.combout(\Add0~45_combout ),
	.cout(\Add0~46 ));
// synopsys translate_off
defparam \Add0~45 .lut_mask = 16'h9617;
defparam \Add0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N0
cycloneive_lcell_comb \Add0~47 (
// Equation(s):
// \Add0~47_combout  = ((Mux24 $ (\Add0~23_combout  $ (!\Add0~46 )))) # (GND)
// \Add0~48  = CARRY((Mux24 & ((\Add0~23_combout ) # (!\Add0~46 ))) # (!Mux24 & (\Add0~23_combout  & !\Add0~46 )))

	.dataa(Mux24),
	.datab(\Add0~23_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~46 ),
	.combout(\Add0~47_combout ),
	.cout(\Add0~48 ));
// synopsys translate_off
defparam \Add0~47 .lut_mask = 16'h698E;
defparam \Add0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N2
cycloneive_lcell_comb \Add0~49 (
// Equation(s):
// \Add0~49_combout  = (\Add0~22_combout  & ((Mux23 & (\Add0~48  & VCC)) # (!Mux23 & (!\Add0~48 )))) # (!\Add0~22_combout  & ((Mux23 & (!\Add0~48 )) # (!Mux23 & ((\Add0~48 ) # (GND)))))
// \Add0~50  = CARRY((\Add0~22_combout  & (!Mux23 & !\Add0~48 )) # (!\Add0~22_combout  & ((!\Add0~48 ) # (!Mux23))))

	.dataa(\Add0~22_combout ),
	.datab(Mux23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~48 ),
	.combout(\Add0~49_combout ),
	.cout(\Add0~50 ));
// synopsys translate_off
defparam \Add0~49 .lut_mask = 16'h9617;
defparam \Add0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N4
cycloneive_lcell_comb \Add0~51 (
// Equation(s):
// \Add0~51_combout  = ((\Add0~21_combout  $ (Mux22 $ (!\Add0~50 )))) # (GND)
// \Add0~52  = CARRY((\Add0~21_combout  & ((Mux22) # (!\Add0~50 ))) # (!\Add0~21_combout  & (Mux22 & !\Add0~50 )))

	.dataa(\Add0~21_combout ),
	.datab(Mux22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~50 ),
	.combout(\Add0~51_combout ),
	.cout(\Add0~52 ));
// synopsys translate_off
defparam \Add0~51 .lut_mask = 16'h698E;
defparam \Add0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N6
cycloneive_lcell_comb \Add0~53 (
// Equation(s):
// \Add0~53_combout  = (Mux21 & ((\Add0~20_combout  & (\Add0~52  & VCC)) # (!\Add0~20_combout  & (!\Add0~52 )))) # (!Mux21 & ((\Add0~20_combout  & (!\Add0~52 )) # (!\Add0~20_combout  & ((\Add0~52 ) # (GND)))))
// \Add0~54  = CARRY((Mux21 & (!\Add0~20_combout  & !\Add0~52 )) # (!Mux21 & ((!\Add0~52 ) # (!\Add0~20_combout ))))

	.dataa(Mux21),
	.datab(\Add0~20_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~52 ),
	.combout(\Add0~53_combout ),
	.cout(\Add0~54 ));
// synopsys translate_off
defparam \Add0~53 .lut_mask = 16'h9617;
defparam \Add0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N8
cycloneive_lcell_comb \Add0~55 (
// Equation(s):
// \Add0~55_combout  = ((Mux20 $ (\Add0~19_combout  $ (!\Add0~54 )))) # (GND)
// \Add0~56  = CARRY((Mux20 & ((\Add0~19_combout ) # (!\Add0~54 ))) # (!Mux20 & (\Add0~19_combout  & !\Add0~54 )))

	.dataa(Mux20),
	.datab(\Add0~19_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~54 ),
	.combout(\Add0~55_combout ),
	.cout(\Add0~56 ));
// synopsys translate_off
defparam \Add0~55 .lut_mask = 16'h698E;
defparam \Add0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N10
cycloneive_lcell_comb \Add0~57 (
// Equation(s):
// \Add0~57_combout  = (\Add0~18_combout  & ((Mux19 & (\Add0~56  & VCC)) # (!Mux19 & (!\Add0~56 )))) # (!\Add0~18_combout  & ((Mux19 & (!\Add0~56 )) # (!Mux19 & ((\Add0~56 ) # (GND)))))
// \Add0~58  = CARRY((\Add0~18_combout  & (!Mux19 & !\Add0~56 )) # (!\Add0~18_combout  & ((!\Add0~56 ) # (!Mux19))))

	.dataa(\Add0~18_combout ),
	.datab(Mux19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~56 ),
	.combout(\Add0~57_combout ),
	.cout(\Add0~58 ));
// synopsys translate_off
defparam \Add0~57 .lut_mask = 16'h9617;
defparam \Add0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N12
cycloneive_lcell_comb \Add0~59 (
// Equation(s):
// \Add0~59_combout  = ((Mux18 $ (\Add0~17_combout  $ (!\Add0~58 )))) # (GND)
// \Add0~60  = CARRY((Mux18 & ((\Add0~17_combout ) # (!\Add0~58 ))) # (!Mux18 & (\Add0~17_combout  & !\Add0~58 )))

	.dataa(Mux18),
	.datab(\Add0~17_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~58 ),
	.combout(\Add0~59_combout ),
	.cout(\Add0~60 ));
// synopsys translate_off
defparam \Add0~59 .lut_mask = 16'h698E;
defparam \Add0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N14
cycloneive_lcell_comb \Add0~61 (
// Equation(s):
// \Add0~61_combout  = (Mux17 & ((\Add0~16_combout  & (\Add0~60  & VCC)) # (!\Add0~16_combout  & (!\Add0~60 )))) # (!Mux17 & ((\Add0~16_combout  & (!\Add0~60 )) # (!\Add0~16_combout  & ((\Add0~60 ) # (GND)))))
// \Add0~62  = CARRY((Mux17 & (!\Add0~16_combout  & !\Add0~60 )) # (!Mux17 & ((!\Add0~60 ) # (!\Add0~16_combout ))))

	.dataa(Mux17),
	.datab(\Add0~16_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~60 ),
	.combout(\Add0~61_combout ),
	.cout(\Add0~62 ));
// synopsys translate_off
defparam \Add0~61 .lut_mask = 16'h9617;
defparam \Add0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N16
cycloneive_lcell_comb \Add0~63 (
// Equation(s):
// \Add0~63_combout  = ((Mux16 $ (\Add0~15_combout  $ (!\Add0~62 )))) # (GND)
// \Add0~64  = CARRY((Mux16 & ((\Add0~15_combout ) # (!\Add0~62 ))) # (!Mux16 & (\Add0~15_combout  & !\Add0~62 )))

	.dataa(Mux16),
	.datab(\Add0~15_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~62 ),
	.combout(\Add0~63_combout ),
	.cout(\Add0~64 ));
// synopsys translate_off
defparam \Add0~63 .lut_mask = 16'h698E;
defparam \Add0~63 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N18
cycloneive_lcell_comb \Add0~65 (
// Equation(s):
// \Add0~65_combout  = (\Add0~14_combout  & ((Mux15 & (\Add0~64  & VCC)) # (!Mux15 & (!\Add0~64 )))) # (!\Add0~14_combout  & ((Mux15 & (!\Add0~64 )) # (!Mux15 & ((\Add0~64 ) # (GND)))))
// \Add0~66  = CARRY((\Add0~14_combout  & (!Mux15 & !\Add0~64 )) # (!\Add0~14_combout  & ((!\Add0~64 ) # (!Mux15))))

	.dataa(\Add0~14_combout ),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~64 ),
	.combout(\Add0~65_combout ),
	.cout(\Add0~66 ));
// synopsys translate_off
defparam \Add0~65 .lut_mask = 16'h9617;
defparam \Add0~65 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N20
cycloneive_lcell_comb \Add0~67 (
// Equation(s):
// \Add0~67_combout  = ((Mux14 $ (\Add0~13_combout  $ (!\Add0~66 )))) # (GND)
// \Add0~68  = CARRY((Mux14 & ((\Add0~13_combout ) # (!\Add0~66 ))) # (!Mux14 & (\Add0~13_combout  & !\Add0~66 )))

	.dataa(Mux14),
	.datab(\Add0~13_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~66 ),
	.combout(\Add0~67_combout ),
	.cout(\Add0~68 ));
// synopsys translate_off
defparam \Add0~67 .lut_mask = 16'h698E;
defparam \Add0~67 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N22
cycloneive_lcell_comb \Add0~69 (
// Equation(s):
// \Add0~69_combout  = (\Add0~12_combout  & ((Mux13 & (\Add0~68  & VCC)) # (!Mux13 & (!\Add0~68 )))) # (!\Add0~12_combout  & ((Mux13 & (!\Add0~68 )) # (!Mux13 & ((\Add0~68 ) # (GND)))))
// \Add0~70  = CARRY((\Add0~12_combout  & (!Mux13 & !\Add0~68 )) # (!\Add0~12_combout  & ((!\Add0~68 ) # (!Mux13))))

	.dataa(\Add0~12_combout ),
	.datab(Mux13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~68 ),
	.combout(\Add0~69_combout ),
	.cout(\Add0~70 ));
// synopsys translate_off
defparam \Add0~69 .lut_mask = 16'h9617;
defparam \Add0~69 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N24
cycloneive_lcell_comb \Add0~71 (
// Equation(s):
// \Add0~71_combout  = ((\Add0~11_combout  $ (Mux12 $ (!\Add0~70 )))) # (GND)
// \Add0~72  = CARRY((\Add0~11_combout  & ((Mux12) # (!\Add0~70 ))) # (!\Add0~11_combout  & (Mux12 & !\Add0~70 )))

	.dataa(\Add0~11_combout ),
	.datab(Mux12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~70 ),
	.combout(\Add0~71_combout ),
	.cout(\Add0~72 ));
// synopsys translate_off
defparam \Add0~71 .lut_mask = 16'h698E;
defparam \Add0~71 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N26
cycloneive_lcell_comb \Add0~73 (
// Equation(s):
// \Add0~73_combout  = (\Add0~10_combout  & ((Mux11 & (\Add0~72  & VCC)) # (!Mux11 & (!\Add0~72 )))) # (!\Add0~10_combout  & ((Mux11 & (!\Add0~72 )) # (!Mux11 & ((\Add0~72 ) # (GND)))))
// \Add0~74  = CARRY((\Add0~10_combout  & (!Mux11 & !\Add0~72 )) # (!\Add0~10_combout  & ((!\Add0~72 ) # (!Mux11))))

	.dataa(\Add0~10_combout ),
	.datab(Mux11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~72 ),
	.combout(\Add0~73_combout ),
	.cout(\Add0~74 ));
// synopsys translate_off
defparam \Add0~73 .lut_mask = 16'h9617;
defparam \Add0~73 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N28
cycloneive_lcell_comb \Add0~75 (
// Equation(s):
// \Add0~75_combout  = ((\Add0~9_combout  $ (Mux10 $ (!\Add0~74 )))) # (GND)
// \Add0~76  = CARRY((\Add0~9_combout  & ((Mux10) # (!\Add0~74 ))) # (!\Add0~9_combout  & (Mux10 & !\Add0~74 )))

	.dataa(\Add0~9_combout ),
	.datab(Mux10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~74 ),
	.combout(\Add0~75_combout ),
	.cout(\Add0~76 ));
// synopsys translate_off
defparam \Add0~75 .lut_mask = 16'h698E;
defparam \Add0~75 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N30
cycloneive_lcell_comb \Add0~77 (
// Equation(s):
// \Add0~77_combout  = (\Add0~8_combout  & ((Mux9 & (\Add0~76  & VCC)) # (!Mux9 & (!\Add0~76 )))) # (!\Add0~8_combout  & ((Mux9 & (!\Add0~76 )) # (!Mux9 & ((\Add0~76 ) # (GND)))))
// \Add0~78  = CARRY((\Add0~8_combout  & (!Mux9 & !\Add0~76 )) # (!\Add0~8_combout  & ((!\Add0~76 ) # (!Mux9))))

	.dataa(\Add0~8_combout ),
	.datab(Mux9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~76 ),
	.combout(\Add0~77_combout ),
	.cout(\Add0~78 ));
// synopsys translate_off
defparam \Add0~77 .lut_mask = 16'h9617;
defparam \Add0~77 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N0
cycloneive_lcell_comb \Add0~79 (
// Equation(s):
// \Add0~79_combout  = ((\Add0~7_combout  $ (Mux8 $ (!\Add0~78 )))) # (GND)
// \Add0~80  = CARRY((\Add0~7_combout  & ((Mux8) # (!\Add0~78 ))) # (!\Add0~7_combout  & (Mux8 & !\Add0~78 )))

	.dataa(\Add0~7_combout ),
	.datab(Mux8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~78 ),
	.combout(\Add0~79_combout ),
	.cout(\Add0~80 ));
// synopsys translate_off
defparam \Add0~79 .lut_mask = 16'h698E;
defparam \Add0~79 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N2
cycloneive_lcell_comb \Add0~81 (
// Equation(s):
// \Add0~81_combout  = (Mux7 & ((\Add0~6_combout  & (\Add0~80  & VCC)) # (!\Add0~6_combout  & (!\Add0~80 )))) # (!Mux7 & ((\Add0~6_combout  & (!\Add0~80 )) # (!\Add0~6_combout  & ((\Add0~80 ) # (GND)))))
// \Add0~82  = CARRY((Mux7 & (!\Add0~6_combout  & !\Add0~80 )) # (!Mux7 & ((!\Add0~80 ) # (!\Add0~6_combout ))))

	.dataa(Mux7),
	.datab(\Add0~6_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~80 ),
	.combout(\Add0~81_combout ),
	.cout(\Add0~82 ));
// synopsys translate_off
defparam \Add0~81 .lut_mask = 16'h9617;
defparam \Add0~81 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N4
cycloneive_lcell_comb \Add0~83 (
// Equation(s):
// \Add0~83_combout  = ((\Add0~5_combout  $ (Mux6 $ (!\Add0~82 )))) # (GND)
// \Add0~84  = CARRY((\Add0~5_combout  & ((Mux6) # (!\Add0~82 ))) # (!\Add0~5_combout  & (Mux6 & !\Add0~82 )))

	.dataa(\Add0~5_combout ),
	.datab(Mux6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~82 ),
	.combout(\Add0~83_combout ),
	.cout(\Add0~84 ));
// synopsys translate_off
defparam \Add0~83 .lut_mask = 16'h698E;
defparam \Add0~83 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N6
cycloneive_lcell_comb \Add0~85 (
// Equation(s):
// \Add0~85_combout  = (Mux5 & ((\Add0~4_combout  & (\Add0~84  & VCC)) # (!\Add0~4_combout  & (!\Add0~84 )))) # (!Mux5 & ((\Add0~4_combout  & (!\Add0~84 )) # (!\Add0~4_combout  & ((\Add0~84 ) # (GND)))))
// \Add0~86  = CARRY((Mux5 & (!\Add0~4_combout  & !\Add0~84 )) # (!Mux5 & ((!\Add0~84 ) # (!\Add0~4_combout ))))

	.dataa(Mux5),
	.datab(\Add0~4_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~84 ),
	.combout(\Add0~85_combout ),
	.cout(\Add0~86 ));
// synopsys translate_off
defparam \Add0~85 .lut_mask = 16'h9617;
defparam \Add0~85 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N8
cycloneive_lcell_comb \Add0~87 (
// Equation(s):
// \Add0~87_combout  = ((\Add0~3_combout  $ (Mux4 $ (!\Add0~86 )))) # (GND)
// \Add0~88  = CARRY((\Add0~3_combout  & ((Mux4) # (!\Add0~86 ))) # (!\Add0~3_combout  & (Mux4 & !\Add0~86 )))

	.dataa(\Add0~3_combout ),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~86 ),
	.combout(\Add0~87_combout ),
	.cout(\Add0~88 ));
// synopsys translate_off
defparam \Add0~87 .lut_mask = 16'h698E;
defparam \Add0~87 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N10
cycloneive_lcell_comb \Add0~89 (
// Equation(s):
// \Add0~89_combout  = (\Add0~2_combout  & ((Mux3 & (\Add0~88  & VCC)) # (!Mux3 & (!\Add0~88 )))) # (!\Add0~2_combout  & ((Mux3 & (!\Add0~88 )) # (!Mux3 & ((\Add0~88 ) # (GND)))))
// \Add0~90  = CARRY((\Add0~2_combout  & (!Mux3 & !\Add0~88 )) # (!\Add0~2_combout  & ((!\Add0~88 ) # (!Mux3))))

	.dataa(\Add0~2_combout ),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~88 ),
	.combout(\Add0~89_combout ),
	.cout(\Add0~90 ));
// synopsys translate_off
defparam \Add0~89 .lut_mask = 16'h9617;
defparam \Add0~89 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N12
cycloneive_lcell_comb \Add0~91 (
// Equation(s):
// \Add0~91_combout  = ((\Add0~1_combout  $ (Mux2 $ (!\Add0~90 )))) # (GND)
// \Add0~92  = CARRY((\Add0~1_combout  & ((Mux2) # (!\Add0~90 ))) # (!\Add0~1_combout  & (Mux2 & !\Add0~90 )))

	.dataa(\Add0~1_combout ),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~90 ),
	.combout(\Add0~91_combout ),
	.cout(\Add0~92 ));
// synopsys translate_off
defparam \Add0~91 .lut_mask = 16'h698E;
defparam \Add0~91 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N14
cycloneive_lcell_comb \Add0~93 (
// Equation(s):
// \Add0~93_combout  = (\Add0~0_combout  & ((Mux1 & (\Add0~92  & VCC)) # (!Mux1 & (!\Add0~92 )))) # (!\Add0~0_combout  & ((Mux1 & (!\Add0~92 )) # (!Mux1 & ((\Add0~92 ) # (GND)))))
// \Add0~94  = CARRY((\Add0~0_combout  & (!Mux1 & !\Add0~92 )) # (!\Add0~0_combout  & ((!\Add0~92 ) # (!Mux1))))

	.dataa(\Add0~0_combout ),
	.datab(Mux1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~92 ),
	.combout(\Add0~93_combout ),
	.cout(\Add0~94 ));
// synopsys translate_off
defparam \Add0~93 .lut_mask = 16'h9617;
defparam \Add0~93 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N10
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (!\Selector99~2_combout  & !\Selector98~2_combout )

	.dataa(Selector991),
	.datab(Selector981),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'h1111;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N20
cycloneive_lcell_comb \ShiftLeft0~38 (
// Equation(s):
// \ShiftLeft0~38_combout  = (\Selector100~4_combout  & ((Mux3))) # (!\Selector100~4_combout  & (Mux2))

	.dataa(Mux2),
	.datab(gnd),
	.datac(Selector1002),
	.datad(Mux3),
	.cin(gnd),
	.combout(\ShiftLeft0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~38 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N24
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (\Mux0~2_combout  & (((!\Mux0~3_combout )))) # (!\Mux0~2_combout  & ((\Mux0~3_combout  & (Mux0)) # (!\Mux0~3_combout  & ((\ShiftLeft0~38_combout )))))

	.dataa(Mux0),
	.datab(\Mux0~2_combout ),
	.datac(\Mux0~3_combout ),
	.datad(\ShiftLeft0~38_combout ),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'h2F2C;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N22
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// \Mux0~9_combout  = (\Mux0~8_combout  & ((\ShiftLeft0~41_combout ) # ((!\Mux0~2_combout )))) # (!\Mux0~8_combout  & (((Mux1 & \Mux0~2_combout ))))

	.dataa(\ShiftLeft0~41_combout ),
	.datab(\Mux0~8_combout ),
	.datac(Mux1),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hB8CC;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N8
cycloneive_lcell_comb \ShiftLeft0~35 (
// Equation(s):
// \ShiftLeft0~35_combout  = (\Selector99~2_combout  & ((Mux10))) # (!\Selector99~2_combout  & (Mux8))

	.dataa(Mux8),
	.datab(Mux10),
	.datac(gnd),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftLeft0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~35 .lut_mask = 16'hCCAA;
defparam \ShiftLeft0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N28
cycloneive_lcell_comb \ShiftLeft0~36 (
// Equation(s):
// \ShiftLeft0~36_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~4_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~35_combout ))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftLeft0~35_combout ),
	.datad(\ShiftLeft0~4_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~36 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N24
cycloneive_lcell_comb \ShiftLeft0~33 (
// Equation(s):
// \ShiftLeft0~33_combout  = (\Selector99~2_combout  & (Mux14)) # (!\Selector99~2_combout  & ((Mux12)))

	.dataa(Selector991),
	.datab(gnd),
	.datac(Mux14),
	.datad(Mux12),
	.cin(gnd),
	.combout(\ShiftLeft0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~33 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N26
cycloneive_lcell_comb \ShiftLeft0~34 (
// Equation(s):
// \ShiftLeft0~34_combout  = (\Selector100~4_combout  & (\ShiftLeft0~1_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~33_combout )))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftLeft0~1_combout ),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~34 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N30
cycloneive_lcell_comb \ShiftLeft0~37 (
// Equation(s):
// \ShiftLeft0~37_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~34_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~36_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~36_combout ),
	.datac(Selector981),
	.datad(\ShiftLeft0~34_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~37 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N16
cycloneive_lcell_comb \ShiftRight0~7 (
// Equation(s):
// \ShiftRight0~7_combout  = (\Mux0~3_combout  & (!\Selector100~4_combout  & (Mux0 & !\Selector97~2_combout )))

	.dataa(\Mux0~3_combout ),
	.datab(Selector1002),
	.datac(Mux0),
	.datad(Selector971),
	.cin(gnd),
	.combout(\ShiftRight0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~7 .lut_mask = 16'h0020;
defparam \ShiftRight0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N30
cycloneive_lcell_comb \ShiftLeft0~42 (
// Equation(s):
// \ShiftLeft0~42_combout  = (!\Selector99~2_combout  & ((\Selector100~4_combout  & (Mux29)) # (!\Selector100~4_combout  & ((Mux28)))))

	.dataa(Selector1002),
	.datab(Selector991),
	.datac(Mux29),
	.datad(Mux28),
	.cin(gnd),
	.combout(\ShiftLeft0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~42 .lut_mask = 16'h3120;
defparam \ShiftLeft0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N24
cycloneive_lcell_comb \ShiftLeft0~43 (
// Equation(s):
// \ShiftLeft0~43_combout  = (\Selector100~4_combout  & (Mux31)) # (!\Selector100~4_combout  & ((Mux30)))

	.dataa(Mux31),
	.datab(gnd),
	.datac(Selector1002),
	.datad(Mux30),
	.cin(gnd),
	.combout(\ShiftLeft0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~43 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N22
cycloneive_lcell_comb \ShiftLeft0~44 (
// Equation(s):
// \ShiftLeft0~44_combout  = (\ShiftLeft0~42_combout ) # ((\Selector99~2_combout  & \ShiftLeft0~43_combout ))

	.dataa(Selector991),
	.datab(gnd),
	.datac(\ShiftLeft0~42_combout ),
	.datad(\ShiftLeft0~43_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~44 .lut_mask = 16'hFAF0;
defparam \ShiftLeft0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N20
cycloneive_lcell_comb \ShiftLeft0~45 (
// Equation(s):
// \ShiftLeft0~45_combout  = (\Selector99~2_combout  & ((Mux26))) # (!\Selector99~2_combout  & (Mux24))

	.dataa(gnd),
	.datab(Mux24),
	.datac(Selector991),
	.datad(Mux26),
	.cin(gnd),
	.combout(\ShiftLeft0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~45 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N18
cycloneive_lcell_comb \ShiftLeft0~46 (
// Equation(s):
// \ShiftLeft0~46_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~22_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~45_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~45_combout ),
	.datac(Selector1002),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~46 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N8
cycloneive_lcell_comb \ShiftLeft0~47 (
// Equation(s):
// \ShiftLeft0~47_combout  = (\Selector98~2_combout  & (\ShiftLeft0~44_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~46_combout )))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~44_combout ),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~47 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N2
cycloneive_lcell_comb \ShiftLeft0~48 (
// Equation(s):
// \ShiftLeft0~48_combout  = (\Selector99~2_combout  & (Mux22)) # (!\Selector99~2_combout  & ((Mux20)))

	.dataa(gnd),
	.datab(Mux22),
	.datac(Mux20),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftLeft0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~48 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N4
cycloneive_lcell_comb \ShiftLeft0~49 (
// Equation(s):
// \ShiftLeft0~49_combout  = (\Selector100~4_combout  & (\ShiftLeft0~26_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~48_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftLeft0~26_combout ),
	.datad(\ShiftLeft0~48_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~49 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N24
cycloneive_lcell_comb \ShiftLeft0~50 (
// Equation(s):
// \ShiftLeft0~50_combout  = (\Selector99~2_combout  & ((Mux18))) # (!\Selector99~2_combout  & (Mux16))

	.dataa(Mux16),
	.datab(gnd),
	.datac(Selector991),
	.datad(Mux18),
	.cin(gnd),
	.combout(\ShiftLeft0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~50 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N10
cycloneive_lcell_comb \ShiftLeft0~51 (
// Equation(s):
// \ShiftLeft0~51_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~29_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~50_combout ))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftLeft0~50_combout ),
	.datad(\ShiftLeft0~29_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~51 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N28
cycloneive_lcell_comb \ShiftLeft0~52 (
// Equation(s):
// \ShiftLeft0~52_combout  = (\Selector98~2_combout  & (\ShiftLeft0~49_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~51_combout )))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~49_combout ),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~52 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N16
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (!\ShiftLeft0~32_combout  & ((\Selector97~2_combout  & (\ShiftLeft0~47_combout )) # (!\Selector97~2_combout  & ((\ShiftLeft0~52_combout )))))

	.dataa(Selector971),
	.datab(\ShiftLeft0~32_combout ),
	.datac(\ShiftLeft0~47_combout ),
	.datad(\ShiftLeft0~52_combout ),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'h3120;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N6
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (\Mux0~7_combout  & (\ShiftRight0~7_combout  & (\Mux0~6_combout ))) # (!\Mux0~7_combout  & (((\Mux0~10_combout ) # (!\Mux0~6_combout ))))

	.dataa(\Mux0~7_combout ),
	.datab(\ShiftRight0~7_combout ),
	.datac(\Mux0~6_combout ),
	.datad(\Mux0~10_combout ),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hD585;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N8
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (\Mux0~5_combout  & (((\Mux0~11_combout )))) # (!\Mux0~5_combout  & ((\Mux0~11_combout  & (\Mux0~9_combout )) # (!\Mux0~11_combout  & ((\ShiftLeft0~37_combout )))))

	.dataa(\Mux0~9_combout ),
	.datab(\Mux0~5_combout ),
	.datac(\ShiftLeft0~37_combout ),
	.datad(\Mux0~11_combout ),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hEE30;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N16
cycloneive_lcell_comb \Add0~95 (
// Equation(s):
// \Add0~95_combout  = Selector3 $ (((\Selector69~0_combout ) # ((Mux321 & \Selector95~0_combout ))))

	.dataa(Selector3),
	.datab(Selector69),
	.datac(Mux32),
	.datad(Selector95),
	.cin(gnd),
	.combout(\Add0~95_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~95 .lut_mask = 16'h5666;
defparam \Add0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N16
cycloneive_lcell_comb \Add0~96 (
// Equation(s):
// \Add0~96_combout  = Mux0 $ (\Add0~94  $ (!\Add0~95_combout ))

	.dataa(Mux0),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add0~95_combout ),
	.cin(\Add0~94 ),
	.combout(\Add0~96_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~96 .lut_mask = 16'h5AA5;
defparam \Add0~96 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N22
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (!Selector1 & (!Selector2 & ((!\ShiftLeft0~32_combout ) # (!Selector3))))

	.dataa(Selector3),
	.datab(Selector1),
	.datac(Selector2),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'h0103;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N6
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (Selector3 & (Selector2 $ (((Mux24) # (\Selector93~1_combout ))))) # (!Selector3 & ((Mux24 & (Selector2 $ (\Selector93~1_combout ))) # (!Mux24 & (Selector2 & \Selector93~1_combout ))))

	.dataa(Selector3),
	.datab(Mux24),
	.datac(Selector2),
	.datad(Selector931),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'h1E68;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N16
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (!Selector2 & !Selector1)

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector2),
	.datad(Selector1),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'h000F;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N22
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (Selector1) # ((Selector3 & !Selector2))

	.dataa(gnd),
	.datab(Selector3),
	.datac(Selector1),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hF0FC;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N24
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (\Mux30~0_combout  & (((!\Mux6~11_combout )))) # (!\Mux30~0_combout  & ((\Mux6~11_combout  & (\Mux24~7_combout )) # (!\Mux6~11_combout  & ((\Add0~47_combout )))))

	.dataa(\Mux24~7_combout ),
	.datab(\Mux30~0_combout ),
	.datac(\Mux6~11_combout ),
	.datad(\Add0~47_combout ),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'h2F2C;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N30
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (!\Selector97~2_combout  & (\Mux0~4_combout  & \ShiftLeft0~47_combout ))

	.dataa(Selector971),
	.datab(gnd),
	.datac(\Mux0~4_combout ),
	.datad(\ShiftLeft0~47_combout ),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'h5000;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N24
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (\Selector97~1_combout ) # ((\Selector96~2_combout ) # ((Mux60 & \Selector100~0_combout )))

	.dataa(Mux60),
	.datab(Selector97),
	.datac(Selector100),
	.datad(Selector961),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hFFEC;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N22
cycloneive_lcell_comb \ShiftRight0~16 (
// Equation(s):
// \ShiftRight0~16_combout  = (\Selector99~2_combout  & ((Mux18))) # (!\Selector99~2_combout  & (Mux20))

	.dataa(Mux20),
	.datab(gnd),
	.datac(Mux18),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftRight0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~16 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N0
cycloneive_lcell_comb \ShiftRight0~15 (
// Equation(s):
// \ShiftRight0~15_combout  = (\Selector99~2_combout  & ((Mux17))) # (!\Selector99~2_combout  & (Mux19))

	.dataa(Mux19),
	.datab(Selector991),
	.datac(gnd),
	.datad(Mux17),
	.cin(gnd),
	.combout(\ShiftRight0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~15 .lut_mask = 16'hEE22;
defparam \ShiftRight0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N4
cycloneive_lcell_comb \ShiftRight0~17 (
// Equation(s):
// \ShiftRight0~17_combout  = (\Selector100~4_combout  & ((\ShiftRight0~15_combout ))) # (!\Selector100~4_combout  & (\ShiftRight0~16_combout ))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftRight0~16_combout ),
	.datad(\ShiftRight0~15_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~17 .lut_mask = 16'hFA50;
defparam \ShiftRight0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N24
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (\Selector96~2_combout ) # ((\Selector98~2_combout  & !\Selector97~2_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(Selector971),
	.datad(Selector961),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hFF0C;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N2
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (\Mux6~18_combout  & (((\Mux6~10_combout )))) # (!\Mux6~18_combout  & ((\Mux6~10_combout  & ((\ShiftRight0~17_combout ))) # (!\Mux6~10_combout  & (\ShiftRight0~20_combout ))))

	.dataa(\ShiftRight0~20_combout ),
	.datab(\Mux6~18_combout ),
	.datac(\ShiftRight0~17_combout ),
	.datad(\Mux6~10_combout ),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hFC22;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N26
cycloneive_lcell_comb \ShiftRight0~12 (
// Equation(s):
// \ShiftRight0~12_combout  = (\Selector99~2_combout  & ((Mux14))) # (!\Selector99~2_combout  & (Mux16))

	.dataa(gnd),
	.datab(Mux16),
	.datac(Mux14),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftRight0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~12 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N6
cycloneive_lcell_comb \ShiftRight0~11 (
// Equation(s):
// \ShiftRight0~11_combout  = (\Selector99~2_combout  & (Mux13)) # (!\Selector99~2_combout  & ((Mux15)))

	.dataa(gnd),
	.datab(Mux13),
	.datac(Mux15),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftRight0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~11 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N8
cycloneive_lcell_comb \ShiftRight0~13 (
// Equation(s):
// \ShiftRight0~13_combout  = (\Selector100~4_combout  & ((\ShiftRight0~11_combout ))) # (!\Selector100~4_combout  & (\ShiftRight0~12_combout ))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftRight0~12_combout ),
	.datad(\ShiftRight0~11_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~13 .lut_mask = 16'hFA50;
defparam \ShiftRight0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N22
cycloneive_lcell_comb \ShiftRight0~8 (
// Equation(s):
// \ShiftRight0~8_combout  = (\Selector99~2_combout  & (Mux9)) # (!\Selector99~2_combout  & ((Mux11)))

	.dataa(Mux9),
	.datab(gnd),
	.datac(Selector991),
	.datad(Mux11),
	.cin(gnd),
	.combout(\ShiftRight0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~8 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N30
cycloneive_lcell_comb \ShiftRight0~9 (
// Equation(s):
// \ShiftRight0~9_combout  = (\Selector99~2_combout  & (Mux10)) # (!\Selector99~2_combout  & ((Mux12)))

	.dataa(Mux10),
	.datab(gnd),
	.datac(Selector991),
	.datad(Mux12),
	.cin(gnd),
	.combout(\ShiftRight0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~9 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N0
cycloneive_lcell_comb \ShiftRight0~10 (
// Equation(s):
// \ShiftRight0~10_combout  = (\Selector100~4_combout  & (\ShiftRight0~8_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~9_combout )))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftRight0~8_combout ),
	.datad(\ShiftRight0~9_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~10 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N14
cycloneive_lcell_comb \ShiftRight0~14 (
// Equation(s):
// \ShiftRight0~14_combout  = (\Selector98~2_combout  & ((\ShiftRight0~10_combout ))) # (!\Selector98~2_combout  & (\ShiftRight0~13_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftRight0~13_combout ),
	.datad(\ShiftRight0~10_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~14 .lut_mask = 16'hFC30;
defparam \ShiftRight0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N12
cycloneive_lcell_comb \ShiftRight0~21 (
// Equation(s):
// \ShiftRight0~21_combout  = (!\Selector98~2_combout  & (!\Selector99~2_combout  & !\Selector100~4_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(Selector991),
	.datad(Selector1002),
	.cin(gnd),
	.combout(\ShiftRight0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~21 .lut_mask = 16'h0003;
defparam \ShiftRight0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N30
cycloneive_lcell_comb \ShiftRight0~22 (
// Equation(s):
// \ShiftRight0~22_combout  = (\Selector100~4_combout  & ((\Selector99~2_combout  & ((Mux1))) # (!\Selector99~2_combout  & (Mux3))))

	.dataa(Selector1002),
	.datab(Selector991),
	.datac(Mux3),
	.datad(Mux1),
	.cin(gnd),
	.combout(\ShiftRight0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~22 .lut_mask = 16'hA820;
defparam \ShiftRight0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N14
cycloneive_lcell_comb \ShiftRight0~23 (
// Equation(s):
// \ShiftRight0~23_combout  = (\Selector99~2_combout  & (Mux2)) # (!\Selector99~2_combout  & ((Mux4)))

	.dataa(Mux2),
	.datab(gnd),
	.datac(Selector991),
	.datad(Mux4),
	.cin(gnd),
	.combout(\ShiftRight0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~23 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N16
cycloneive_lcell_comb \ShiftRight0~24 (
// Equation(s):
// \ShiftRight0~24_combout  = (\ShiftRight0~22_combout ) # ((!\Selector100~4_combout  & \ShiftRight0~23_combout ))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftRight0~22_combout ),
	.datad(\ShiftRight0~23_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~24 .lut_mask = 16'hF5F0;
defparam \ShiftRight0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N8
cycloneive_lcell_comb \ShiftRight0~25 (
// Equation(s):
// \ShiftRight0~25_combout  = (\Selector99~2_combout  & (Mux5)) # (!\Selector99~2_combout  & ((Mux7)))

	.dataa(gnd),
	.datab(Selector991),
	.datac(Mux5),
	.datad(Mux7),
	.cin(gnd),
	.combout(\ShiftRight0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~25 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N14
cycloneive_lcell_comb \ShiftRight0~26 (
// Equation(s):
// \ShiftRight0~26_combout  = (\Selector99~2_combout  & ((Mux6))) # (!\Selector99~2_combout  & (Mux8))

	.dataa(Mux8),
	.datab(Selector991),
	.datac(gnd),
	.datad(Mux6),
	.cin(gnd),
	.combout(\ShiftRight0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~26 .lut_mask = 16'hEE22;
defparam \ShiftRight0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N20
cycloneive_lcell_comb \ShiftRight0~27 (
// Equation(s):
// \ShiftRight0~27_combout  = (\Selector100~4_combout  & (\ShiftRight0~25_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~26_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftRight0~25_combout ),
	.datad(\ShiftRight0~26_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~27 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N14
cycloneive_lcell_comb \ShiftRight0~28 (
// Equation(s):
// \ShiftRight0~28_combout  = (\Selector98~2_combout  & (\ShiftRight0~24_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~27_combout )))

	.dataa(Selector981),
	.datab(\ShiftRight0~24_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~27_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~28 .lut_mask = 16'hDD88;
defparam \ShiftRight0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N4
cycloneive_lcell_comb \ShiftRight0~29 (
// Equation(s):
// \ShiftRight0~29_combout  = (\Selector97~2_combout  & (Mux0 & (\ShiftRight0~21_combout ))) # (!\Selector97~2_combout  & (((\ShiftRight0~28_combout ))))

	.dataa(Mux0),
	.datab(Selector971),
	.datac(\ShiftRight0~21_combout ),
	.datad(\ShiftRight0~28_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~29 .lut_mask = 16'hB380;
defparam \ShiftRight0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N28
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (\Mux6~18_combout  & ((\Mux24~4_combout  & ((\ShiftRight0~29_combout ))) # (!\Mux24~4_combout  & (\ShiftRight0~14_combout )))) # (!\Mux6~18_combout  & (\Mux24~4_combout ))

	.dataa(\Mux6~18_combout ),
	.datab(\Mux24~4_combout ),
	.datac(\ShiftRight0~14_combout ),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hEC64;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N30
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (\ShiftLeft0~24_combout  & (!\Selector97~2_combout  & \Mux0~4_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~24_combout ),
	.datac(Selector971),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'h0C00;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N28
cycloneive_lcell_comb \ShiftRight0~39 (
// Equation(s):
// \ShiftRight0~39_combout  = (\Selector99~2_combout  & (Mux3)) # (!\Selector99~2_combout  & ((Mux5)))

	.dataa(gnd),
	.datab(Mux3),
	.datac(Selector991),
	.datad(Mux5),
	.cin(gnd),
	.combout(\ShiftRight0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~39 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N26
cycloneive_lcell_comb \ShiftRight0~40 (
// Equation(s):
// \ShiftRight0~40_combout  = (\Selector100~4_combout  & (\ShiftRight0~23_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~39_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~23_combout ),
	.datac(Selector1002),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~40 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N28
cycloneive_lcell_comb \ShiftRight0~41 (
// Equation(s):
// \ShiftRight0~41_combout  = (\Selector99~2_combout  & (Mux7)) # (!\Selector99~2_combout  & ((Mux9)))

	.dataa(gnd),
	.datab(Mux7),
	.datac(Mux9),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftRight0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~41 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N28
cycloneive_lcell_comb \ShiftRight0~42 (
// Equation(s):
// \ShiftRight0~42_combout  = (\Selector100~4_combout  & (\ShiftRight0~26_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~41_combout )))

	.dataa(Selector1002),
	.datab(\ShiftRight0~26_combout ),
	.datac(\ShiftRight0~41_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~42 .lut_mask = 16'hD8D8;
defparam \ShiftRight0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N22
cycloneive_lcell_comb \ShiftRight0~43 (
// Equation(s):
// \ShiftRight0~43_combout  = (\Selector98~2_combout  & (\ShiftRight0~40_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~42_combout )))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftRight0~40_combout ),
	.datad(\ShiftRight0~42_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~43 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N8
cycloneive_lcell_comb \ShiftRight0~44 (
// Equation(s):
// \ShiftRight0~44_combout  = (\Selector97~2_combout  & (\Mux0~3_combout  & ((\ShiftRight0~6_combout )))) # (!\Selector97~2_combout  & (((\ShiftRight0~43_combout ))))

	.dataa(Selector971),
	.datab(\Mux0~3_combout ),
	.datac(\ShiftRight0~43_combout ),
	.datad(\ShiftRight0~6_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~44 .lut_mask = 16'hD850;
defparam \ShiftRight0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N26
cycloneive_lcell_comb \ShiftRight0~30 (
// Equation(s):
// \ShiftRight0~30_combout  = (\Selector99~2_combout  & (Mux19)) # (!\Selector99~2_combout  & ((Mux21)))

	.dataa(Mux19),
	.datab(gnd),
	.datac(Selector991),
	.datad(Mux21),
	.cin(gnd),
	.combout(\ShiftRight0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~30 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N4
cycloneive_lcell_comb \ShiftRight0~31 (
// Equation(s):
// \ShiftRight0~31_combout  = (\Selector100~4_combout  & ((\ShiftRight0~16_combout ))) # (!\Selector100~4_combout  & (\ShiftRight0~30_combout ))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftRight0~30_combout ),
	.datad(\ShiftRight0~16_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~31 .lut_mask = 16'hFC30;
defparam \ShiftRight0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N2
cycloneive_lcell_comb \ShiftRight0~32 (
// Equation(s):
// \ShiftRight0~32_combout  = (\Selector99~2_combout  & (Mux11)) # (!\Selector99~2_combout  & ((Mux13)))

	.dataa(gnd),
	.datab(Mux11),
	.datac(Mux13),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftRight0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~32 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N0
cycloneive_lcell_comb \ShiftRight0~33 (
// Equation(s):
// \ShiftRight0~33_combout  = (\Selector100~4_combout  & (\ShiftRight0~9_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~32_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftRight0~9_combout ),
	.datad(\ShiftRight0~32_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~33 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N18
cycloneive_lcell_comb \ShiftRight0~34 (
// Equation(s):
// \ShiftRight0~34_combout  = (\Selector99~2_combout  & (Mux15)) # (!\Selector99~2_combout  & ((Mux17)))

	.dataa(Mux15),
	.datab(gnd),
	.datac(Selector991),
	.datad(Mux17),
	.cin(gnd),
	.combout(\ShiftRight0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~34 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N12
cycloneive_lcell_comb \ShiftRight0~35 (
// Equation(s):
// \ShiftRight0~35_combout  = (\Selector100~4_combout  & (\ShiftRight0~12_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~34_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftRight0~12_combout ),
	.datad(\ShiftRight0~34_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~35 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N10
cycloneive_lcell_comb \ShiftRight0~36 (
// Equation(s):
// \ShiftRight0~36_combout  = (\Selector98~2_combout  & (\ShiftRight0~33_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~35_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~33_combout ),
	.datac(Selector981),
	.datad(\ShiftRight0~35_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~36 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N18
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (\Mux6~10_combout  & (((\Mux6~18_combout )))) # (!\Mux6~10_combout  & ((\Mux6~18_combout  & ((\ShiftRight0~36_combout ))) # (!\Mux6~18_combout  & (\ShiftRight0~38_combout ))))

	.dataa(\ShiftRight0~38_combout ),
	.datab(\Mux6~10_combout ),
	.datac(\Mux6~18_combout ),
	.datad(\ShiftRight0~36_combout ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hF2C2;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N20
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Mux6~10_combout  & ((\Mux25~0_combout  & (\ShiftRight0~44_combout )) # (!\Mux25~0_combout  & ((\ShiftRight0~31_combout ))))) # (!\Mux6~10_combout  & (((\Mux25~0_combout ))))

	.dataa(\Mux6~10_combout ),
	.datab(\ShiftRight0~44_combout ),
	.datac(\ShiftRight0~31_combout ),
	.datad(\Mux25~0_combout ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hDDA0;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N0
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (\Selector94~1_combout  & (Selector2 $ (((Mux25) # (Selector3))))) # (!\Selector94~1_combout  & ((Selector2 & (Mux25 $ (Selector3))) # (!Selector2 & (Mux25 & Selector3))))

	.dataa(Selector941),
	.datab(Selector2),
	.datac(Mux25),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'h3668;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N2
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (\Mux6~11_combout  & (\Mux25~3_combout  & ((!\Mux30~0_combout )))) # (!\Mux6~11_combout  & (((\Add0~45_combout ) # (\Mux30~0_combout ))))

	.dataa(\Mux6~11_combout ),
	.datab(\Mux25~3_combout ),
	.datac(\Add0~45_combout ),
	.datad(\Mux30~0_combout ),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'h55D8;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N14
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (Selector3 & (Selector2 $ (((Mux26) # (\Selector95~3_combout ))))) # (!Selector3 & ((Mux26 & (Selector2 $ (\Selector95~3_combout ))) # (!Mux26 & (Selector2 & \Selector95~3_combout ))))

	.dataa(Selector3),
	.datab(Mux26),
	.datac(Selector2),
	.datad(Selector952),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'h1E68;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N20
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (\Mux6~11_combout  & (!\Mux30~0_combout  & (\Mux26~3_combout ))) # (!\Mux6~11_combout  & ((\Mux30~0_combout ) # ((\Add0~43_combout ))))

	.dataa(\Mux6~11_combout ),
	.datab(\Mux30~0_combout ),
	.datac(\Mux26~3_combout ),
	.datad(\Add0~43_combout ),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'h7564;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N10
cycloneive_lcell_comb \ShiftLeft0~53 (
// Equation(s):
// \ShiftLeft0~53_combout  = (\Selector99~2_combout  & ((Mux29))) # (!\Selector99~2_combout  & (Mux27))

	.dataa(gnd),
	.datab(Mux27),
	.datac(Selector991),
	.datad(Mux29),
	.cin(gnd),
	.combout(\ShiftLeft0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~53 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N12
cycloneive_lcell_comb \ShiftLeft0~21 (
// Equation(s):
// \ShiftLeft0~21_combout  = (\Selector99~2_combout  & ((Mux28))) # (!\Selector99~2_combout  & (Mux26))

	.dataa(gnd),
	.datab(Selector991),
	.datac(Mux26),
	.datad(Mux28),
	.cin(gnd),
	.combout(\ShiftLeft0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~21 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N0
cycloneive_lcell_comb \ShiftLeft0~54 (
// Equation(s):
// \ShiftLeft0~54_combout  = (\Selector100~4_combout  & (\ShiftLeft0~53_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~21_combout )))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftLeft0~53_combout ),
	.datad(\ShiftLeft0~21_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~54 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N8
cycloneive_lcell_comb \ShiftLeft0~55 (
// Equation(s):
// \ShiftLeft0~55_combout  = (\Selector98~2_combout  & (!\Selector99~2_combout  & (\ShiftLeft0~43_combout ))) # (!\Selector98~2_combout  & (((\ShiftLeft0~54_combout ))))

	.dataa(Selector991),
	.datab(\ShiftLeft0~43_combout ),
	.datac(Selector981),
	.datad(\ShiftLeft0~54_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~55 .lut_mask = 16'h4F40;
defparam \ShiftLeft0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N8
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (!\Selector97~2_combout  & (\Mux0~4_combout  & \ShiftLeft0~55_combout ))

	.dataa(Selector971),
	.datab(gnd),
	.datac(\Mux0~4_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'h5000;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N16
cycloneive_lcell_comb \ShiftRight0~52 (
// Equation(s):
// \ShiftRight0~52_combout  = (\Selector99~2_combout  & ((\Selector100~4_combout  & ((Mux23))) # (!\Selector100~4_combout  & (Mux24))))

	.dataa(Mux24),
	.datab(Selector1002),
	.datac(Mux23),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~52 .lut_mask = 16'hE200;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N6
cycloneive_lcell_comb \ShiftRight0~53 (
// Equation(s):
// \ShiftRight0~53_combout  = (\Selector100~4_combout  & (Mux25)) # (!\Selector100~4_combout  & ((Mux26)))

	.dataa(Mux25),
	.datab(gnd),
	.datac(Selector1002),
	.datad(Mux26),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~53 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N2
cycloneive_lcell_comb \ShiftRight0~54 (
// Equation(s):
// \ShiftRight0~54_combout  = (\ShiftRight0~52_combout ) # ((!\Selector99~2_combout  & \ShiftRight0~53_combout ))

	.dataa(Selector991),
	.datab(gnd),
	.datac(\ShiftRight0~52_combout ),
	.datad(\ShiftRight0~53_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~54 .lut_mask = 16'hF5F0;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N12
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (\Mux6~18_combout  & (((\Mux6~10_combout )))) # (!\Mux6~18_combout  & ((\Mux6~10_combout  & (\ShiftRight0~51_combout )) # (!\Mux6~10_combout  & ((\ShiftRight0~54_combout )))))

	.dataa(\ShiftRight0~51_combout ),
	.datab(\Mux6~18_combout ),
	.datac(\ShiftRight0~54_combout ),
	.datad(\Mux6~10_combout ),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hEE30;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N10
cycloneive_lcell_comb \ShiftRight0~45 (
// Equation(s):
// \ShiftRight0~45_combout  = (\Selector99~2_combout  & ((Mux12))) # (!\Selector99~2_combout  & (Mux14))

	.dataa(Selector991),
	.datab(gnd),
	.datac(Mux14),
	.datad(Mux12),
	.cin(gnd),
	.combout(\ShiftRight0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~45 .lut_mask = 16'hFA50;
defparam \ShiftRight0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N4
cycloneive_lcell_comb \ShiftRight0~46 (
// Equation(s):
// \ShiftRight0~46_combout  = (\Selector100~4_combout  & (\ShiftRight0~32_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~45_combout )))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftRight0~32_combout ),
	.datad(\ShiftRight0~45_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~46 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N6
cycloneive_lcell_comb \ShiftRight0~47 (
// Equation(s):
// \ShiftRight0~47_combout  = (\Selector99~2_combout  & (Mux16)) # (!\Selector99~2_combout  & ((Mux18)))

	.dataa(gnd),
	.datab(Mux16),
	.datac(Mux18),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftRight0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~47 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N28
cycloneive_lcell_comb \ShiftRight0~48 (
// Equation(s):
// \ShiftRight0~48_combout  = (\Selector100~4_combout  & ((\ShiftRight0~34_combout ))) # (!\Selector100~4_combout  & (\ShiftRight0~47_combout ))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftRight0~47_combout ),
	.datad(\ShiftRight0~34_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~48 .lut_mask = 16'hFC30;
defparam \ShiftRight0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N14
cycloneive_lcell_comb \ShiftRight0~49 (
// Equation(s):
// \ShiftRight0~49_combout  = (\Selector98~2_combout  & (\ShiftRight0~46_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~48_combout )))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftRight0~46_combout ),
	.datad(\ShiftRight0~48_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~49 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N22
cycloneive_lcell_comb \ShiftRight0~55 (
// Equation(s):
// \ShiftRight0~55_combout  = (\Selector99~2_combout  & (Mux4)) # (!\Selector99~2_combout  & ((Mux6)))

	.dataa(gnd),
	.datab(Selector991),
	.datac(Mux4),
	.datad(Mux6),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~55 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N24
cycloneive_lcell_comb \ShiftRight0~56 (
// Equation(s):
// \ShiftRight0~56_combout  = (\Selector100~4_combout  & ((\ShiftRight0~39_combout ))) # (!\Selector100~4_combout  & (\ShiftRight0~55_combout ))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftRight0~55_combout ),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~56 .lut_mask = 16'hFC30;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N0
cycloneive_lcell_comb \ShiftRight0~57 (
// Equation(s):
// \ShiftRight0~57_combout  = (\Selector99~2_combout  & (Mux8)) # (!\Selector99~2_combout  & ((Mux10)))

	.dataa(gnd),
	.datab(Selector991),
	.datac(Mux8),
	.datad(Mux10),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~57 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N20
cycloneive_lcell_comb \ShiftRight0~58 (
// Equation(s):
// \ShiftRight0~58_combout  = (\Selector100~4_combout  & ((\ShiftRight0~41_combout ))) # (!\Selector100~4_combout  & (\ShiftRight0~57_combout ))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftRight0~57_combout ),
	.datad(\ShiftRight0~41_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~58 .lut_mask = 16'hFA50;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N8
cycloneive_lcell_comb \ShiftRight0~59 (
// Equation(s):
// \ShiftRight0~59_combout  = (\Selector98~2_combout  & (\ShiftRight0~56_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~58_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~56_combout ),
	.datac(Selector981),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~59 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N18
cycloneive_lcell_comb \ShiftRight0~60 (
// Equation(s):
// \ShiftRight0~60_combout  = (!\Selector100~4_combout  & ((\Selector99~2_combout  & ((Mux0))) # (!\Selector99~2_combout  & (Mux2))))

	.dataa(Mux2),
	.datab(Selector991),
	.datac(Selector1002),
	.datad(Mux0),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~60 .lut_mask = 16'h0E02;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N16
cycloneive_lcell_comb \ShiftRight0~61 (
// Equation(s):
// \ShiftRight0~61_combout  = (\ShiftRight0~60_combout ) # ((!\Selector99~2_combout  & (\Selector100~4_combout  & Mux1)))

	.dataa(Selector991),
	.datab(Selector1002),
	.datac(Mux1),
	.datad(\ShiftRight0~60_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~61 .lut_mask = 16'hFF40;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N10
cycloneive_lcell_comb \ShiftRight0~62 (
// Equation(s):
// \ShiftRight0~62_combout  = (\Selector97~2_combout  & (!\Selector98~2_combout  & ((\ShiftRight0~61_combout )))) # (!\Selector97~2_combout  & (((\ShiftRight0~59_combout ))))

	.dataa(Selector981),
	.datab(Selector971),
	.datac(\ShiftRight0~59_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~62 .lut_mask = 16'h7430;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N10
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (\Mux26~0_combout  & (((\ShiftRight0~62_combout )) # (!\Mux6~18_combout ))) # (!\Mux26~0_combout  & (\Mux6~18_combout  & (\ShiftRight0~49_combout )))

	.dataa(\Mux26~0_combout ),
	.datab(\Mux6~18_combout ),
	.datac(\ShiftRight0~49_combout ),
	.datad(\ShiftRight0~62_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hEA62;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N14
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (Selector3 & (Selector2 $ (((\Selector96~2_combout ) # (Mux27))))) # (!Selector3 & ((Selector2 & (\Selector96~2_combout  $ (Mux27))) # (!Selector2 & (\Selector96~2_combout  & Mux27))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(Selector961),
	.datad(Mux27),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'h5668;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N10
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (\Mux30~0_combout  & (!\Mux6~11_combout )) # (!\Mux30~0_combout  & ((\Mux6~11_combout  & ((\Mux27~3_combout ))) # (!\Mux6~11_combout  & (\Add0~41_combout ))))

	.dataa(\Mux30~0_combout ),
	.datab(\Mux6~11_combout ),
	.datac(\Add0~41_combout ),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'h7632;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N8
cycloneive_lcell_comb \ShiftLeft0~57 (
// Equation(s):
// \ShiftLeft0~57_combout  = (\Selector99~2_combout  & ((Mux30))) # (!\Selector99~2_combout  & (Mux28))

	.dataa(gnd),
	.datab(Mux28),
	.datac(Selector991),
	.datad(Mux30),
	.cin(gnd),
	.combout(\ShiftLeft0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~57 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N14
cycloneive_lcell_comb \ShiftLeft0~58 (
// Equation(s):
// \ShiftLeft0~58_combout  = (\Selector100~4_combout  & (\ShiftLeft0~57_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~53_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftLeft0~57_combout ),
	.datad(\ShiftLeft0~53_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~58 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N16
cycloneive_lcell_comb \ShiftLeft0~56 (
// Equation(s):
// \ShiftLeft0~56_combout  = (\Selector98~2_combout  & (!\Selector99~2_combout  & !\Selector100~4_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(Selector991),
	.datad(Selector1002),
	.cin(gnd),
	.combout(\ShiftLeft0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~56 .lut_mask = 16'h000C;
defparam \ShiftLeft0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N16
cycloneive_lcell_comb \ShiftLeft0~59 (
// Equation(s):
// \ShiftLeft0~59_combout  = (Mux31 & ((\ShiftLeft0~56_combout ) # ((!\Selector98~2_combout  & \ShiftLeft0~58_combout )))) # (!Mux31 & (!\Selector98~2_combout  & (\ShiftLeft0~58_combout )))

	.dataa(Mux31),
	.datab(Selector981),
	.datac(\ShiftLeft0~58_combout ),
	.datad(\ShiftLeft0~56_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~59 .lut_mask = 16'hBA30;
defparam \ShiftLeft0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N28
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (\Mux0~4_combout  & (!\Selector97~2_combout  & \ShiftLeft0~59_combout ))

	.dataa(gnd),
	.datab(\Mux0~4_combout ),
	.datac(Selector971),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'h0C00;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N20
cycloneive_lcell_comb \ShiftRight0~18 (
// Equation(s):
// \ShiftRight0~18_combout  = (\Selector99~2_combout  & ((Mux21))) # (!\Selector99~2_combout  & (Mux23))

	.dataa(Mux23),
	.datab(gnd),
	.datac(Selector991),
	.datad(Mux21),
	.cin(gnd),
	.combout(\ShiftRight0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~18 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N14
cycloneive_lcell_comb \ShiftRight0~63 (
// Equation(s):
// \ShiftRight0~63_combout  = (\Selector100~4_combout  & (\ShiftRight0~50_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~18_combout )))

	.dataa(\ShiftRight0~50_combout ),
	.datab(Selector1002),
	.datac(gnd),
	.datad(\ShiftRight0~18_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~63 .lut_mask = 16'hBB88;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N8
cycloneive_lcell_comb \ShiftRight0~74 (
// Equation(s):
// \ShiftRight0~74_combout  = (\ShiftRight0~73_combout ) # ((\Selector99~2_combout  & \ShiftRight0~6_combout ))

	.dataa(\ShiftRight0~73_combout ),
	.datab(gnd),
	.datac(Selector991),
	.datad(\ShiftRight0~6_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~74 .lut_mask = 16'hFAAA;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N2
cycloneive_lcell_comb \ShiftRight0~71 (
// Equation(s):
// \ShiftRight0~71_combout  = (\Selector100~4_combout  & (\ShiftRight0~57_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~8_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftRight0~57_combout ),
	.datad(\ShiftRight0~8_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~71 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N10
cycloneive_lcell_comb \ShiftRight0~70 (
// Equation(s):
// \ShiftRight0~70_combout  = (\Selector100~4_combout  & (\ShiftRight0~55_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~25_combout )))

	.dataa(\ShiftRight0~55_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~25_combout ),
	.datad(Selector1002),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~70 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N10
cycloneive_lcell_comb \ShiftRight0~72 (
// Equation(s):
// \ShiftRight0~72_combout  = (\Selector98~2_combout  & ((\ShiftRight0~70_combout ))) # (!\Selector98~2_combout  & (\ShiftRight0~71_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftRight0~71_combout ),
	.datad(\ShiftRight0~70_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~72 .lut_mask = 16'hFC30;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N4
cycloneive_lcell_comb \ShiftRight0~75 (
// Equation(s):
// \ShiftRight0~75_combout  = (\Selector97~2_combout  & (!\Selector98~2_combout  & (\ShiftRight0~74_combout ))) # (!\Selector97~2_combout  & (((\ShiftRight0~72_combout ))))

	.dataa(Selector971),
	.datab(Selector981),
	.datac(\ShiftRight0~74_combout ),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~75 .lut_mask = 16'h7520;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N26
cycloneive_lcell_comb \ShiftRight0~64 (
// Equation(s):
// \ShiftRight0~64_combout  = (\Selector100~4_combout  & (\ShiftRight0~45_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~11_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftRight0~45_combout ),
	.datad(\ShiftRight0~11_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~64 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N16
cycloneive_lcell_comb \ShiftRight0~65 (
// Equation(s):
// \ShiftRight0~65_combout  = (\Selector100~4_combout  & (\ShiftRight0~47_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~15_combout )))

	.dataa(\ShiftRight0~47_combout ),
	.datab(gnd),
	.datac(Selector1002),
	.datad(\ShiftRight0~15_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~65 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N18
cycloneive_lcell_comb \ShiftRight0~66 (
// Equation(s):
// \ShiftRight0~66_combout  = (\Selector98~2_combout  & (\ShiftRight0~64_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~65_combout )))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftRight0~64_combout ),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~66 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N12
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (\Mux6~10_combout  & (((\Mux6~18_combout )))) # (!\Mux6~10_combout  & ((\Mux6~18_combout  & ((\ShiftRight0~66_combout ))) # (!\Mux6~18_combout  & (\ShiftRight0~69_combout ))))

	.dataa(\ShiftRight0~69_combout ),
	.datab(\Mux6~10_combout ),
	.datac(\Mux6~18_combout ),
	.datad(\ShiftRight0~66_combout ),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hF2C2;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N2
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (\Mux6~10_combout  & ((\Mux27~0_combout  & ((\ShiftRight0~75_combout ))) # (!\Mux27~0_combout  & (\ShiftRight0~63_combout )))) # (!\Mux6~10_combout  & (((\Mux27~0_combout ))))

	.dataa(\Mux6~10_combout ),
	.datab(\ShiftRight0~63_combout ),
	.datac(\ShiftRight0~75_combout ),
	.datad(\Mux27~0_combout ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hF588;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N30
cycloneive_lcell_comb \Mux6~20 (
// Equation(s):
// \Mux6~20_combout  = (!Selector1 & (!Selector2 & ((\Mux0~4_combout ) # (!Selector3))))

	.dataa(Selector3),
	.datab(Selector1),
	.datac(Selector2),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux6~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~20 .lut_mask = 16'h0301;
defparam \Mux6~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N22
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (Selector3 & (Selector2 $ (((Mux4) # (\Selector73~1_combout ))))) # (!Selector3 & ((Mux4 & (Selector2 $ (\Selector73~1_combout ))) # (!Mux4 & (Selector2 & \Selector73~1_combout ))))

	.dataa(Selector3),
	.datab(Mux4),
	.datac(Selector2),
	.datad(Selector731),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'h1E68;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N24
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (\Mux30~0_combout  & (((!\Mux6~11_combout )))) # (!\Mux30~0_combout  & ((\Mux6~11_combout  & (\Mux4~4_combout )) # (!\Mux6~11_combout  & ((\Add0~87_combout )))))

	.dataa(\Mux4~4_combout ),
	.datab(\Mux30~0_combout ),
	.datac(\Mux6~11_combout ),
	.datad(\Add0~87_combout ),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'h2F2C;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N12
cycloneive_lcell_comb \ShiftRight0~76 (
// Equation(s):
// \ShiftRight0~76_combout  = (\Selector98~2_combout  & (\ShiftLeft0~56_combout  & (Mux0))) # (!\Selector98~2_combout  & ((\ShiftRight0~24_combout ) # ((\ShiftLeft0~56_combout  & Mux0))))

	.dataa(Selector981),
	.datab(\ShiftLeft0~56_combout ),
	.datac(Mux0),
	.datad(\ShiftRight0~24_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~76 .lut_mask = 16'hD5C0;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N22
cycloneive_lcell_comb \ShiftRight0~104 (
// Equation(s):
// \ShiftRight0~104_combout  = (!\Selector97~1_combout  & (\ShiftRight0~76_combout  & ((!\Selector100~0_combout ) # (!Mux60))))

	.dataa(Mux60),
	.datab(Selector97),
	.datac(Selector100),
	.datad(\ShiftRight0~76_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~104 .lut_mask = 16'h1300;
defparam \ShiftRight0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N22
cycloneive_lcell_comb \ShiftLeft0~39 (
// Equation(s):
// \ShiftLeft0~39_combout  = (\Selector99~2_combout  & ((\Selector100~4_combout  & ((Mux7))) # (!\Selector100~4_combout  & (Mux6))))

	.dataa(Selector1002),
	.datab(Mux6),
	.datac(Mux7),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftLeft0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~39 .lut_mask = 16'hE400;
defparam \ShiftLeft0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N24
cycloneive_lcell_comb \ShiftLeft0~40 (
// Equation(s):
// \ShiftLeft0~40_combout  = (\Selector100~4_combout  & (Mux5)) # (!\Selector100~4_combout  & ((Mux4)))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(Mux5),
	.datad(Mux4),
	.cin(gnd),
	.combout(\ShiftLeft0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~40 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N14
cycloneive_lcell_comb \ShiftLeft0~41 (
// Equation(s):
// \ShiftLeft0~41_combout  = (\ShiftLeft0~39_combout ) # ((!\Selector99~2_combout  & \ShiftLeft0~40_combout ))

	.dataa(gnd),
	.datab(Selector991),
	.datac(\ShiftLeft0~39_combout ),
	.datad(\ShiftLeft0~40_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~41 .lut_mask = 16'hF3F0;
defparam \ShiftLeft0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N18
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (\Mux6~18_combout  & (((\Mux6~10_combout )))) # (!\Mux6~18_combout  & ((\Mux6~10_combout  & ((\ShiftLeft0~36_combout ))) # (!\Mux6~10_combout  & (\ShiftLeft0~41_combout ))))

	.dataa(\Mux6~18_combout ),
	.datab(\ShiftLeft0~41_combout ),
	.datac(\Mux6~10_combout ),
	.datad(\ShiftLeft0~36_combout ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hF4A4;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N22
cycloneive_lcell_comb \ShiftLeft0~60 (
// Equation(s):
// \ShiftLeft0~60_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~51_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~34_combout ))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~34_combout ),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~60 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N0
cycloneive_lcell_comb \ShiftLeft0~61 (
// Equation(s):
// \ShiftLeft0~61_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~46_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~49_combout ))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~49_combout ),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~61 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N6
cycloneive_lcell_comb \ShiftLeft0~62 (
// Equation(s):
// \ShiftLeft0~62_combout  = (\Selector97~2_combout  & (!\Selector98~2_combout  & (\ShiftLeft0~44_combout ))) # (!\Selector97~2_combout  & (((\ShiftLeft0~61_combout ))))

	.dataa(Selector981),
	.datab(Selector971),
	.datac(\ShiftLeft0~44_combout ),
	.datad(\ShiftLeft0~61_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~62 .lut_mask = 16'h7340;
defparam \ShiftLeft0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N12
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (\Mux6~18_combout  & ((\Mux4~2_combout  & ((\ShiftLeft0~62_combout ))) # (!\Mux4~2_combout  & (\ShiftLeft0~60_combout )))) # (!\Mux6~18_combout  & (\Mux4~2_combout ))

	.dataa(\Mux6~18_combout ),
	.datab(\Mux4~2_combout ),
	.datac(\ShiftLeft0~60_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hEC64;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N2
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (!\ShiftLeft0~18_combout  & (!\ShiftLeft0~15_combout  & (!\ShiftLeft0~16_combout  & \Mux4~3_combout )))

	.dataa(\ShiftLeft0~18_combout ),
	.datab(\ShiftLeft0~15_combout ),
	.datac(\ShiftLeft0~16_combout ),
	.datad(\Mux4~3_combout ),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'h0100;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N30
cycloneive_lcell_comb \ShiftLeft0~64 (
// Equation(s):
// \ShiftLeft0~64_combout  = (\Selector98~2_combout  & (\ShiftLeft0~23_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~27_combout )))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~23_combout ),
	.datad(\ShiftLeft0~27_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~64 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N30
cycloneive_lcell_comb \ShiftLeft0~65 (
// Equation(s):
// \ShiftLeft0~65_combout  = (\Selector97~2_combout  & (!\Selector98~2_combout  & (\ShiftLeft0~20_combout ))) # (!\Selector97~2_combout  & (((\ShiftLeft0~64_combout ))))

	.dataa(Selector971),
	.datab(Selector981),
	.datac(\ShiftLeft0~20_combout ),
	.datad(\ShiftLeft0~64_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~65 .lut_mask = 16'h7520;
defparam \ShiftLeft0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N4
cycloneive_lcell_comb \ShiftLeft0~63 (
// Equation(s):
// \ShiftLeft0~63_combout  = (\Selector98~2_combout  & (\ShiftLeft0~30_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~2_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~30_combout ),
	.datac(Selector981),
	.datad(\ShiftLeft0~2_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~63 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N22
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (\Mux6~10_combout  & (\Mux6~18_combout )) # (!\Mux6~10_combout  & ((\Mux6~18_combout  & (\ShiftLeft0~63_combout )) # (!\Mux6~18_combout  & ((\ShiftLeft0~10_combout )))))

	.dataa(\Mux6~10_combout ),
	.datab(\Mux6~18_combout ),
	.datac(\ShiftLeft0~63_combout ),
	.datad(\ShiftLeft0~10_combout ),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hD9C8;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N16
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (\Mux6~10_combout  & ((\Mux5~2_combout  & ((\ShiftLeft0~65_combout ))) # (!\Mux5~2_combout  & (\ShiftLeft0~5_combout )))) # (!\Mux6~10_combout  & (((\Mux5~2_combout ))))

	.dataa(\Mux6~10_combout ),
	.datab(\ShiftLeft0~5_combout ),
	.datac(\ShiftLeft0~65_combout ),
	.datad(\Mux5~2_combout ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hF588;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N18
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (!\ShiftLeft0~18_combout  & (!\ShiftLeft0~16_combout  & (!\ShiftLeft0~15_combout  & \Mux5~3_combout )))

	.dataa(\ShiftLeft0~18_combout ),
	.datab(\ShiftLeft0~16_combout ),
	.datac(\ShiftLeft0~15_combout ),
	.datad(\Mux5~3_combout ),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'h0100;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N2
cycloneive_lcell_comb \ShiftRight0~77 (
// Equation(s):
// \ShiftRight0~77_combout  = (\Selector98~2_combout  & (((!\Selector99~2_combout  & \ShiftRight0~6_combout )))) # (!\Selector98~2_combout  & (\ShiftRight0~40_combout ))

	.dataa(\ShiftRight0~40_combout ),
	.datab(Selector981),
	.datac(Selector991),
	.datad(\ShiftRight0~6_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~77 .lut_mask = 16'h2E22;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N10
cycloneive_lcell_comb \ShiftRight0~105 (
// Equation(s):
// \ShiftRight0~105_combout  = (!\Selector97~1_combout  & (\ShiftRight0~77_combout  & ((!\Selector100~0_combout ) # (!Mux60))))

	.dataa(Mux60),
	.datab(Selector100),
	.datac(Selector97),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~105 .lut_mask = 16'h0700;
defparam \ShiftRight0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N20
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (Mux5 & (Selector2 $ (((Selector3) # (\Selector74~1_combout ))))) # (!Mux5 & ((Selector2 & (Selector3 $ (\Selector74~1_combout ))) # (!Selector2 & (Selector3 & \Selector74~1_combout ))))

	.dataa(Mux5),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector741),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'h3668;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N26
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (\Mux6~11_combout  & (\Mux5~4_combout  & (!\Mux30~0_combout ))) # (!\Mux6~11_combout  & (((\Mux30~0_combout ) # (\Add0~85_combout ))))

	.dataa(\Mux6~11_combout ),
	.datab(\Mux5~4_combout ),
	.datac(\Mux30~0_combout ),
	.datad(\Add0~85_combout ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'h5D58;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N20
cycloneive_lcell_comb \ShiftRight0~78 (
// Equation(s):
// \ShiftRight0~78_combout  = (!\Selector97~2_combout  & ((\Selector98~2_combout  & (\ShiftRight0~61_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~56_combout )))))

	.dataa(Selector981),
	.datab(\ShiftRight0~61_combout ),
	.datac(Selector971),
	.datad(\ShiftRight0~56_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~78 .lut_mask = 16'h0D08;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N16
cycloneive_lcell_comb \ShiftLeft0~68 (
// Equation(s):
// \ShiftLeft0~68_combout  = (\Selector99~2_combout  & ((Mux17))) # (!\Selector99~2_combout  & (Mux15))

	.dataa(Selector991),
	.datab(gnd),
	.datac(Mux15),
	.datad(Mux17),
	.cin(gnd),
	.combout(\ShiftLeft0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~68 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N0
cycloneive_lcell_comb \ShiftLeft0~69 (
// Equation(s):
// \ShiftLeft0~69_combout  = (\Selector100~4_combout  & (\ShiftLeft0~68_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~0_combout )))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftLeft0~68_combout ),
	.datad(\ShiftLeft0~0_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~69 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N6
cycloneive_lcell_comb \ShiftLeft0~28 (
// Equation(s):
// \ShiftLeft0~28_combout  = (\Selector99~2_combout  & (Mux20)) # (!\Selector99~2_combout  & ((Mux18)))

	.dataa(Selector991),
	.datab(gnd),
	.datac(Mux20),
	.datad(Mux18),
	.cin(gnd),
	.combout(\ShiftLeft0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~28 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N6
cycloneive_lcell_comb \ShiftLeft0~66 (
// Equation(s):
// \ShiftLeft0~66_combout  = (\Selector99~2_combout  & (Mux21)) # (!\Selector99~2_combout  & ((Mux19)))

	.dataa(Mux21),
	.datab(gnd),
	.datac(Mux19),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftLeft0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~66 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N2
cycloneive_lcell_comb \ShiftLeft0~67 (
// Equation(s):
// \ShiftLeft0~67_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~66_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~28_combout ))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftLeft0~28_combout ),
	.datad(\ShiftLeft0~66_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~67 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N20
cycloneive_lcell_comb \ShiftLeft0~70 (
// Equation(s):
// \ShiftLeft0~70_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~67_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~69_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftLeft0~69_combout ),
	.datad(\ShiftLeft0~67_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~70 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N2
cycloneive_lcell_comb \ShiftLeft0~73 (
// Equation(s):
// \ShiftLeft0~73_combout  = (!\Selector100~4_combout  & ((\Selector99~2_combout  & (Mux8)) # (!\Selector99~2_combout  & ((Mux6)))))

	.dataa(Selector991),
	.datab(Mux8),
	.datac(Selector1002),
	.datad(Mux6),
	.cin(gnd),
	.combout(\ShiftLeft0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~73 .lut_mask = 16'h0D08;
defparam \ShiftLeft0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N0
cycloneive_lcell_comb \ShiftLeft0~75 (
// Equation(s):
// \ShiftLeft0~75_combout  = (\ShiftLeft0~73_combout ) # ((\ShiftLeft0~74_combout  & \Selector100~4_combout ))

	.dataa(\ShiftLeft0~74_combout ),
	.datab(gnd),
	.datac(Selector1002),
	.datad(\ShiftLeft0~73_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~75 .lut_mask = 16'hFFA0;
defparam \ShiftLeft0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N12
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (\Mux6~10_combout  & ((\ShiftLeft0~72_combout ) # ((\Mux6~18_combout )))) # (!\Mux6~10_combout  & (((!\Mux6~18_combout  & \ShiftLeft0~75_combout ))))

	.dataa(\ShiftLeft0~72_combout ),
	.datab(\Mux6~10_combout ),
	.datac(\Mux6~18_combout ),
	.datad(\ShiftLeft0~75_combout ),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hCBC8;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N24
cycloneive_lcell_comb \ShiftLeft0~76 (
// Equation(s):
// \ShiftLeft0~76_combout  = (\Selector99~2_combout  & ((Mux25))) # (!\Selector99~2_combout  & (Mux23))

	.dataa(Mux23),
	.datab(gnd),
	.datac(Mux25),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftLeft0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~76 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N12
cycloneive_lcell_comb \ShiftLeft0~77 (
// Equation(s):
// \ShiftLeft0~77_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~76_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~25_combout ))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftLeft0~25_combout ),
	.datad(\ShiftLeft0~76_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~77 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N6
cycloneive_lcell_comb \ShiftLeft0~78 (
// Equation(s):
// \ShiftLeft0~78_combout  = (\Selector98~2_combout  & (\ShiftLeft0~54_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~77_combout )))

	.dataa(Selector981),
	.datab(\ShiftLeft0~54_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~77_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~78 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N28
cycloneive_lcell_comb \ShiftLeft0~79 (
// Equation(s):
// \ShiftLeft0~79_combout  = (\Selector97~2_combout  & (\Mux0~3_combout  & (\ShiftLeft0~43_combout ))) # (!\Selector97~2_combout  & (((\ShiftLeft0~78_combout ))))

	.dataa(Selector971),
	.datab(\Mux0~3_combout ),
	.datac(\ShiftLeft0~43_combout ),
	.datad(\ShiftLeft0~78_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~79 .lut_mask = 16'hD580;
defparam \ShiftLeft0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N18
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (\Mux6~18_combout  & ((\Mux6~12_combout  & ((\ShiftLeft0~79_combout ))) # (!\Mux6~12_combout  & (\ShiftLeft0~70_combout )))) # (!\Mux6~18_combout  & (((\Mux6~12_combout ))))

	.dataa(\Mux6~18_combout ),
	.datab(\ShiftLeft0~70_combout ),
	.datac(\Mux6~12_combout ),
	.datad(\ShiftLeft0~79_combout ),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hF858;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N8
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// \Mux6~19_combout  = (!\ShiftLeft0~16_combout  & (!\ShiftLeft0~15_combout  & (!\ShiftLeft0~18_combout  & \Mux6~13_combout )))

	.dataa(\ShiftLeft0~16_combout ),
	.datab(\ShiftLeft0~15_combout ),
	.datac(\ShiftLeft0~18_combout ),
	.datad(\Mux6~13_combout ),
	.cin(gnd),
	.combout(\Mux6~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'h0100;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N28
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (\Selector75~1_combout  & (Selector2 $ (((Selector3) # (Mux6))))) # (!\Selector75~1_combout  & ((Selector3 & (Selector2 $ (Mux6))) # (!Selector3 & (Selector2 & Mux6))))

	.dataa(Selector751),
	.datab(Selector3),
	.datac(Selector2),
	.datad(Mux6),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'h1E68;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N18
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (\Mux30~0_combout  & (((!\Mux6~11_combout )))) # (!\Mux30~0_combout  & ((\Mux6~11_combout  & ((\Mux6~14_combout ))) # (!\Mux6~11_combout  & (\Add0~83_combout ))))

	.dataa(\Mux30~0_combout ),
	.datab(\Add0~83_combout ),
	.datac(\Mux6~11_combout ),
	.datad(\Mux6~14_combout ),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'h5E0E;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N14
cycloneive_lcell_comb \ShiftRight0~79 (
// Equation(s):
// \ShiftRight0~79_combout  = (!\Selector97~2_combout  & ((\Selector98~2_combout  & (\ShiftRight0~74_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~70_combout )))))

	.dataa(Selector971),
	.datab(\ShiftRight0~74_combout ),
	.datac(Selector981),
	.datad(\ShiftRight0~70_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~79 .lut_mask = 16'h4540;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N16
cycloneive_lcell_comb \ShiftLeft0~85 (
// Equation(s):
// \ShiftLeft0~85_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~45_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~76_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~76_combout ),
	.datac(Selector1002),
	.datad(\ShiftLeft0~45_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~85 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N28
cycloneive_lcell_comb \ShiftLeft0~86 (
// Equation(s):
// \ShiftLeft0~86_combout  = (\Selector98~2_combout  & (\ShiftLeft0~58_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~85_combout )))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftLeft0~58_combout ),
	.datad(\ShiftLeft0~85_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~86 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N6
cycloneive_lcell_comb \ShiftLeft0~87 (
// Equation(s):
// \ShiftLeft0~87_combout  = (\Selector97~2_combout  & (\ShiftRight0~21_combout  & (Mux31))) # (!\Selector97~2_combout  & (((\ShiftLeft0~86_combout ))))

	.dataa(\ShiftRight0~21_combout ),
	.datab(Mux31),
	.datac(Selector971),
	.datad(\ShiftLeft0~86_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~87 .lut_mask = 16'h8F80;
defparam \ShiftLeft0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N12
cycloneive_lcell_comb \ShiftLeft0~74 (
// Equation(s):
// \ShiftLeft0~74_combout  = (\Selector99~2_combout  & ((Mux9))) # (!\Selector99~2_combout  & (Mux7))

	.dataa(gnd),
	.datab(Mux7),
	.datac(Mux9),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftLeft0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~74 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N14
cycloneive_lcell_comb \ShiftLeft0~84 (
// Equation(s):
// \ShiftLeft0~84_combout  = (\Selector100~4_combout  & (\ShiftLeft0~35_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~74_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftLeft0~35_combout ),
	.datad(\ShiftLeft0~74_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~84 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N30
cycloneive_lcell_comb \ShiftLeft0~81 (
// Equation(s):
// \ShiftLeft0~81_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~48_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~66_combout ))

	.dataa(\ShiftLeft0~66_combout ),
	.datab(Selector1002),
	.datac(gnd),
	.datad(\ShiftLeft0~48_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~81 .lut_mask = 16'hEE22;
defparam \ShiftLeft0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N12
cycloneive_lcell_comb \ShiftLeft0~82 (
// Equation(s):
// \ShiftLeft0~82_combout  = (\Selector100~4_combout  & ((\ShiftLeft0~50_combout ))) # (!\Selector100~4_combout  & (\ShiftLeft0~68_combout ))

	.dataa(\ShiftLeft0~68_combout ),
	.datab(Selector1002),
	.datac(gnd),
	.datad(\ShiftLeft0~50_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~82 .lut_mask = 16'hEE22;
defparam \ShiftLeft0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N30
cycloneive_lcell_comb \ShiftLeft0~83 (
// Equation(s):
// \ShiftLeft0~83_combout  = (\Selector98~2_combout  & (\ShiftLeft0~81_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~82_combout )))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftLeft0~81_combout ),
	.datad(\ShiftLeft0~82_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~83 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N20
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (\Mux6~18_combout  & ((\Mux6~10_combout ) # ((\ShiftLeft0~83_combout )))) # (!\Mux6~18_combout  & (!\Mux6~10_combout  & (\ShiftLeft0~84_combout )))

	.dataa(\Mux6~18_combout ),
	.datab(\Mux6~10_combout ),
	.datac(\ShiftLeft0~84_combout ),
	.datad(\ShiftLeft0~83_combout ),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hBA98;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N18
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (\Mux6~10_combout  & ((\Mux7~2_combout  & ((\ShiftLeft0~87_combout ))) # (!\Mux7~2_combout  & (\ShiftLeft0~80_combout )))) # (!\Mux6~10_combout  & (((\Mux7~2_combout ))))

	.dataa(\ShiftLeft0~80_combout ),
	.datab(\Mux6~10_combout ),
	.datac(\ShiftLeft0~87_combout ),
	.datad(\Mux7~2_combout ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hF388;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N0
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (!\ShiftLeft0~18_combout  & (!\ShiftLeft0~15_combout  & (!\ShiftLeft0~16_combout  & \Mux7~3_combout )))

	.dataa(\ShiftLeft0~18_combout ),
	.datab(\ShiftLeft0~15_combout ),
	.datac(\ShiftLeft0~16_combout ),
	.datad(\Mux7~3_combout ),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'h0100;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N4
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (Selector3 & (Selector2 $ (((\Selector76~1_combout ) # (Mux7))))) # (!Selector3 & ((\Selector76~1_combout  & (Mux7 $ (Selector2))) # (!\Selector76~1_combout  & (Mux7 & Selector2))))

	.dataa(Selector3),
	.datab(Selector761),
	.datac(Mux7),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'h16E8;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N22
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (\Mux30~0_combout  & (!\Mux6~11_combout )) # (!\Mux30~0_combout  & ((\Mux6~11_combout  & (\Mux7~4_combout )) # (!\Mux6~11_combout  & ((\Add0~81_combout )))))

	.dataa(\Mux30~0_combout ),
	.datab(\Mux6~11_combout ),
	.datac(\Mux7~4_combout ),
	.datad(\Add0~81_combout ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'h7362;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N22
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (Mux271) # ((Mux251) # ((Mux261) # (Mux241)))

	.dataa(Mux271),
	.datab(Mux251),
	.datac(Mux261),
	.datad(Mux241),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'hFFFE;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N10
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// \Equal0~1_combout  = (Mux64) # ((Mux71) # ((Mux410) # (Mux510)))

	.dataa(Mux64),
	.datab(Mux71),
	.datac(Mux410),
	.datad(Mux510),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'hFFFE;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N20
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (Mux3 & (Selector2 $ (((Selector3) # (\Selector72~1_combout ))))) # (!Mux3 & ((Selector3 & (Selector2 $ (\Selector72~1_combout ))) # (!Selector3 & (Selector2 & \Selector72~1_combout ))))

	.dataa(Mux3),
	.datab(Selector3),
	.datac(Selector2),
	.datad(Selector721),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'h1E68;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N6
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (Selector3) # (Selector2)

	.dataa(Selector3),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hFFAA;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N10
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (!Selector0 & (!Selector1 & ((\Mux2~0_combout ) # (!\ShiftLeft0~32_combout ))))

	.dataa(\Mux2~0_combout ),
	.datab(Selector0),
	.datac(Selector1),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'h0203;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N14
cycloneive_lcell_comb \ShiftLeft0~88 (
// Equation(s):
// \ShiftLeft0~88_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~85_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~81_combout ))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~81_combout ),
	.datad(\ShiftLeft0~85_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~88 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N14
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (\Selector97~2_combout  & ((\ShiftLeft0~59_combout ))) # (!\Selector97~2_combout  & (\ShiftLeft0~88_combout ))

	.dataa(Selector971),
	.datab(gnd),
	.datac(\ShiftLeft0~88_combout ),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hFA50;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N6
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (\Selector97~2_combout ) # ((!\Selector98~2_combout  & \Selector99~2_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(Selector991),
	.datad(Selector971),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hFF30;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N30
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (\Selector97~1_combout ) # ((\Selector98~2_combout ) # ((Mux60 & \Selector100~0_combout )))

	.dataa(Mux60),
	.datab(Selector97),
	.datac(Selector100),
	.datad(Selector981),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hFFEC;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N2
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (\Mux2~1_combout  & (((!\Mux2~2_combout )))) # (!\Mux2~1_combout  & ((\Mux2~2_combout  & ((\ShiftLeft0~84_combout ))) # (!\Mux2~2_combout  & (\ShiftLeft0~7_combout ))))

	.dataa(\ShiftLeft0~7_combout ),
	.datab(\ShiftLeft0~84_combout ),
	.datac(\Mux2~1_combout ),
	.datad(\Mux2~2_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'h0CFA;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N16
cycloneive_lcell_comb \ShiftLeft0~89 (
// Equation(s):
// \ShiftLeft0~89_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~82_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~80_combout ))

	.dataa(\ShiftLeft0~80_combout ),
	.datab(Selector981),
	.datac(\ShiftLeft0~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~89 .lut_mask = 16'hE2E2;
defparam \ShiftLeft0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N14
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (\Mux2~1_combout  & ((\Mux3~1_combout  & (\ShiftLeft0~9_combout )) # (!\Mux3~1_combout  & ((\ShiftLeft0~89_combout ))))) # (!\Mux2~1_combout  & (((\Mux3~1_combout ))))

	.dataa(\ShiftLeft0~9_combout ),
	.datab(\Mux2~1_combout ),
	.datac(\Mux3~1_combout ),
	.datad(\ShiftLeft0~89_combout ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hBCB0;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N6
cycloneive_lcell_comb \ShiftRight0~73 (
// Equation(s):
// \ShiftRight0~73_combout  = (!\Selector99~2_combout  & ((\Selector100~4_combout  & (Mux2)) # (!\Selector100~4_combout  & ((Mux3)))))

	.dataa(Mux2),
	.datab(Mux3),
	.datac(Selector1002),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~73 .lut_mask = 16'h00AC;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N16
cycloneive_lcell_comb \ShiftRight0~80 (
// Equation(s):
// \ShiftRight0~80_combout  = (!\Mux2~2_combout  & ((\ShiftRight0~73_combout ) # ((\Selector99~2_combout  & \ShiftRight0~6_combout ))))

	.dataa(Selector991),
	.datab(\Mux2~2_combout ),
	.datac(\ShiftRight0~6_combout ),
	.datad(\ShiftRight0~73_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~80 .lut_mask = 16'h3320;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N10
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (Selector2) # ((Selector3 & \Mux0~4_combout ))

	.dataa(Selector3),
	.datab(gnd),
	.datac(Selector2),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hFAF0;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N24
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (\Mux2~4_combout  & (((\Add0~89_combout ) # (!\Mux2~3_combout )))) # (!\Mux2~4_combout  & (\ShiftRight0~80_combout  & (\Mux2~3_combout )))

	.dataa(\Mux2~4_combout ),
	.datab(\ShiftRight0~80_combout ),
	.datac(\Mux2~3_combout ),
	.datad(\Add0~89_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hEA4A;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N2
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (\Mux2~0_combout  & (((\Mux3~3_combout )))) # (!\Mux2~0_combout  & ((\Mux3~3_combout  & (\Mux3~0_combout )) # (!\Mux3~3_combout  & ((\Mux3~2_combout )))))

	.dataa(\Mux2~0_combout ),
	.datab(\Mux3~0_combout ),
	.datac(\Mux3~2_combout ),
	.datad(\Mux3~3_combout ),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hEE50;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N10
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (Mux2 & (Selector2 $ (((Selector3) # (\Selector71~1_combout ))))) # (!Mux2 & ((Selector2 & (Selector3 $ (\Selector71~1_combout ))) # (!Selector2 & (Selector3 & \Selector71~1_combout ))))

	.dataa(Mux2),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector711),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'h3668;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N24
cycloneive_lcell_comb \ShiftLeft0~90 (
// Equation(s):
// \ShiftLeft0~90_combout  = (\Selector98~2_combout  & ((\ShiftLeft0~77_combout ))) # (!\Selector98~2_combout  & (\ShiftLeft0~67_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~67_combout ),
	.datac(Selector981),
	.datad(\ShiftLeft0~77_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~90 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N8
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (\Selector97~2_combout  & ((\ShiftLeft0~55_combout ))) # (!\Selector97~2_combout  & (\ShiftLeft0~90_combout ))

	.dataa(gnd),
	.datab(Selector971),
	.datac(\ShiftLeft0~90_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hFC30;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N8
cycloneive_lcell_comb \ShiftLeft0~71 (
// Equation(s):
// \ShiftLeft0~71_combout  = (\Selector99~2_combout  & (Mux13)) # (!\Selector99~2_combout  & ((Mux11)))

	.dataa(Mux13),
	.datab(gnd),
	.datac(Mux11),
	.datad(Selector991),
	.cin(gnd),
	.combout(\ShiftLeft0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~71 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N6
cycloneive_lcell_comb \ShiftLeft0~72 (
// Equation(s):
// \ShiftLeft0~72_combout  = (\Selector100~4_combout  & (\ShiftLeft0~71_combout )) # (!\Selector100~4_combout  & ((\ShiftLeft0~3_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftLeft0~71_combout ),
	.datad(\ShiftLeft0~3_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~72 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N24
cycloneive_lcell_comb \ShiftLeft0~91 (
// Equation(s):
// \ShiftLeft0~91_combout  = (\Selector98~2_combout  & (\ShiftLeft0~69_combout )) # (!\Selector98~2_combout  & ((\ShiftLeft0~72_combout )))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftLeft0~69_combout ),
	.datad(\ShiftLeft0~72_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~91 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N26
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (\Mux2~6_combout  & ((\ShiftLeft0~40_combout ) # ((!\Mux2~1_combout )))) # (!\Mux2~6_combout  & (((\Mux2~1_combout  & \ShiftLeft0~91_combout ))))

	.dataa(\Mux2~6_combout ),
	.datab(\ShiftLeft0~40_combout ),
	.datac(\Mux2~1_combout ),
	.datad(\ShiftLeft0~91_combout ),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hDA8A;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N20
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (Selector2) # ((\Selector96~2_combout  & !Selector3))

	.dataa(Selector2),
	.datab(Selector961),
	.datac(gnd),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hAAEE;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N0
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (\Mux2~4_combout  & (((\Add0~91_combout ) # (!\Mux2~3_combout )))) # (!\Mux2~4_combout  & (\ShiftRight0~81_combout  & (\Mux2~3_combout )))

	.dataa(\ShiftRight0~81_combout ),
	.datab(\Mux2~4_combout ),
	.datac(\Mux2~3_combout ),
	.datad(\Add0~91_combout ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hEC2C;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N18
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// \Mux2~9_combout  = (\Mux2~0_combout  & (((\Mux2~8_combout )))) # (!\Mux2~0_combout  & ((\Mux2~8_combout  & (\Mux2~5_combout )) # (!\Mux2~8_combout  & ((\Mux2~7_combout )))))

	.dataa(\Mux2~0_combout ),
	.datab(\Mux2~5_combout ),
	.datac(\Mux2~7_combout ),
	.datad(\Mux2~8_combout ),
	.cin(gnd),
	.combout(\Mux2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hEE50;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N26
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = Selector3 $ (((\Selector92~0_combout ) # ((\Selector95~0_combout  & Mux55))))

	.dataa(Selector95),
	.datab(Selector3),
	.datac(Mux55),
	.datad(Selector92),
	.cin(gnd),
	.combout(\Add0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h336C;
defparam \Add0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N20
cycloneive_lcell_comb \ShiftRight0~82 (
// Equation(s):
// \ShiftRight0~82_combout  = (\Selector98~2_combout  & (\ShiftRight0~71_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~64_combout )))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftRight0~71_combout ),
	.datad(\ShiftRight0~64_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~82 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N16
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (!Selector3) # (!\Mux0~4_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux0~4_combout ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'h0FFF;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N8
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = ((!\Mux0~4_combout  & !\ShiftLeft0~32_combout )) # (!Selector3)

	.dataa(gnd),
	.datab(Selector3),
	.datac(\Mux0~4_combout ),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'h333F;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N18
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (\Mux0~4_combout  & \ShiftLeft0~87_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux0~4_combout ),
	.datad(\ShiftLeft0~87_combout ),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hF000;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N30
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (\Mux18~4_combout  & (\Mux18~3_combout  & (\ShiftRight0~79_combout ))) # (!\Mux18~4_combout  & (((\Mux23~4_combout )) # (!\Mux18~3_combout )))

	.dataa(\Mux18~4_combout ),
	.datab(\Mux18~3_combout ),
	.datac(\ShiftRight0~79_combout ),
	.datad(\Mux23~4_combout ),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hD591;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N24
cycloneive_lcell_comb \ShiftRight0~83 (
// Equation(s):
// \ShiftRight0~83_combout  = (\Selector98~2_combout  & ((\ShiftRight0~65_combout ))) # (!\Selector98~2_combout  & (\ShiftRight0~63_combout ))

	.dataa(Selector981),
	.datab(\ShiftRight0~63_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~83 .lut_mask = 16'hEE44;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N20
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (\Mux18~2_combout  & (((\Mux23~5_combout )))) # (!\Mux18~2_combout  & ((\Mux23~5_combout  & ((\ShiftRight0~83_combout ))) # (!\Mux23~5_combout  & (\ShiftRight0~82_combout ))))

	.dataa(\ShiftRight0~82_combout ),
	.datab(\Mux18~2_combout ),
	.datac(\Mux23~5_combout ),
	.datad(\ShiftRight0~83_combout ),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hF2C2;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N4
cycloneive_lcell_comb \Add0~21 (
// Equation(s):
// \Add0~21_combout  = Selector3 $ (((\Selector91~0_combout ) # ((Mux54 & \Selector95~0_combout ))))

	.dataa(Selector3),
	.datab(Mux54),
	.datac(Selector91),
	.datad(Selector95),
	.cin(gnd),
	.combout(\Add0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~21 .lut_mask = 16'h565A;
defparam \Add0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N6
cycloneive_lcell_comb \ShiftRight0~50 (
// Equation(s):
// \ShiftRight0~50_combout  = (\Selector99~2_combout  & (Mux20)) # (!\Selector99~2_combout  & ((Mux22)))

	.dataa(Mux20),
	.datab(gnd),
	.datac(Selector991),
	.datad(Mux22),
	.cin(gnd),
	.combout(\ShiftRight0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~50 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N16
cycloneive_lcell_comb \ShiftRight0~51 (
// Equation(s):
// \ShiftRight0~51_combout  = (\Selector100~4_combout  & (\ShiftRight0~30_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~50_combout )))

	.dataa(gnd),
	.datab(Selector1002),
	.datac(\ShiftRight0~30_combout ),
	.datad(\ShiftRight0~50_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~51 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N8
cycloneive_lcell_comb \ShiftRight0~85 (
// Equation(s):
// \ShiftRight0~85_combout  = (\Selector98~2_combout  & ((\ShiftRight0~48_combout ))) # (!\Selector98~2_combout  & (\ShiftRight0~51_combout ))

	.dataa(Selector981),
	.datab(\ShiftRight0~51_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~48_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~85 .lut_mask = 16'hEE44;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N10
cycloneive_lcell_comb \ShiftRight0~84 (
// Equation(s):
// \ShiftRight0~84_combout  = (\Selector98~2_combout  & ((\ShiftRight0~58_combout ))) # (!\Selector98~2_combout  & (\ShiftRight0~46_combout ))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftRight0~46_combout ),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~84 .lut_mask = 16'hFA50;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N26
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (Selector3 & ((\Selector97~2_combout ) # ((\Selector96~2_combout ) # (\ShiftLeft0~32_combout ))))

	.dataa(Selector971),
	.datab(Selector3),
	.datac(Selector961),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hCCC8;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N12
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (\Mux0~4_combout  & \ShiftLeft0~79_combout )

	.dataa(\Mux0~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ShiftLeft0~79_combout ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hAA00;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N6
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (\Mux18~3_combout  & ((\Mux18~4_combout  & (\ShiftRight0~78_combout )) # (!\Mux18~4_combout  & ((\Mux22~2_combout ))))) # (!\Mux18~3_combout  & (((!\Mux18~4_combout ))))

	.dataa(\ShiftRight0~78_combout ),
	.datab(\Mux18~3_combout ),
	.datac(\Mux18~4_combout ),
	.datad(\Mux22~2_combout ),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'h8F83;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N20
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (\Mux18~2_combout  & (((\Mux22~3_combout )))) # (!\Mux18~2_combout  & ((\Mux22~3_combout  & (\ShiftRight0~85_combout )) # (!\Mux22~3_combout  & ((\ShiftRight0~84_combout )))))

	.dataa(\ShiftRight0~85_combout ),
	.datab(\ShiftRight0~84_combout ),
	.datac(\Mux18~2_combout ),
	.datad(\Mux22~3_combout ),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hFA0C;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N22
cycloneive_lcell_comb \ShiftRight0~87 (
// Equation(s):
// \ShiftRight0~87_combout  = (\Selector98~2_combout  & ((\ShiftRight0~35_combout ))) # (!\Selector98~2_combout  & (\ShiftRight0~31_combout ))

	.dataa(Selector981),
	.datab(gnd),
	.datac(\ShiftRight0~31_combout ),
	.datad(\ShiftRight0~35_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~87 .lut_mask = 16'hFA50;
defparam \ShiftRight0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N6
cycloneive_lcell_comb \ShiftRight0~86 (
// Equation(s):
// \ShiftRight0~86_combout  = (\Selector98~2_combout  & ((\ShiftRight0~42_combout ))) # (!\Selector98~2_combout  & (\ShiftRight0~33_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftRight0~33_combout ),
	.datad(\ShiftRight0~42_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~86 .lut_mask = 16'hFC30;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N24
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (\ShiftLeft0~65_combout  & \Mux0~4_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~65_combout ),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hF000;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N2
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (\Mux18~3_combout  & ((\Mux18~4_combout  & (\ShiftRight0~105_combout )) # (!\Mux18~4_combout  & ((\Mux21~2_combout ))))) # (!\Mux18~3_combout  & (((!\Mux18~4_combout ))))

	.dataa(\ShiftRight0~105_combout ),
	.datab(\Mux18~3_combout ),
	.datac(\Mux18~4_combout ),
	.datad(\Mux21~2_combout ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'h8F83;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N4
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (\Mux18~2_combout  & (((\Mux21~3_combout )))) # (!\Mux18~2_combout  & ((\Mux21~3_combout  & (\ShiftRight0~87_combout )) # (!\Mux21~3_combout  & ((\ShiftRight0~86_combout )))))

	.dataa(\ShiftRight0~87_combout ),
	.datab(\Mux18~2_combout ),
	.datac(\ShiftRight0~86_combout ),
	.datad(\Mux21~3_combout ),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hEE30;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N30
cycloneive_lcell_comb \ShiftRight0~89 (
// Equation(s):
// \ShiftRight0~89_combout  = (\Selector98~2_combout  & (\ShiftRight0~13_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~17_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~13_combout ),
	.datac(\ShiftRight0~17_combout ),
	.datad(Selector981),
	.cin(gnd),
	.combout(\ShiftRight0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~89 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N4
cycloneive_lcell_comb \ShiftRight0~88 (
// Equation(s):
// \ShiftRight0~88_combout  = (\Selector98~2_combout  & ((\ShiftRight0~27_combout ))) # (!\Selector98~2_combout  & (\ShiftRight0~10_combout ))

	.dataa(Selector981),
	.datab(\ShiftRight0~10_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~27_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~88 .lut_mask = 16'hEE44;
defparam \ShiftRight0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N18
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (\Mux0~4_combout  & \ShiftLeft0~62_combout )

	.dataa(\Mux0~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hAA00;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N24
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (\Mux18~3_combout  & ((\Mux18~4_combout  & (\ShiftRight0~104_combout )) # (!\Mux18~4_combout  & ((\Mux20~2_combout ))))) # (!\Mux18~3_combout  & (((!\Mux18~4_combout ))))

	.dataa(\ShiftRight0~104_combout ),
	.datab(\Mux18~3_combout ),
	.datac(\Mux18~4_combout ),
	.datad(\Mux20~2_combout ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'h8F83;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N2
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (\Mux18~2_combout  & (((\Mux20~3_combout )))) # (!\Mux18~2_combout  & ((\Mux20~3_combout  & (\ShiftRight0~89_combout )) # (!\Mux20~3_combout  & ((\ShiftRight0~88_combout )))))

	.dataa(\ShiftRight0~89_combout ),
	.datab(\ShiftRight0~88_combout ),
	.datac(\Mux18~2_combout ),
	.datad(\Mux20~3_combout ),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hFA0C;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N16
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = Selector3 $ (((\Selector88~0_combout ) # ((Mux51 & \Selector95~0_combout ))))

	.dataa(Selector3),
	.datab(Mux51),
	.datac(Selector88),
	.datad(Selector95),
	.cin(gnd),
	.combout(\Add0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h565A;
defparam \Add0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N4
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (\Mux18~4_combout  & (((\ShiftRight0~80_combout  & \Mux18~3_combout )))) # (!\Mux18~4_combout  & ((\Mux19~2_combout ) # ((!\Mux18~3_combout ))))

	.dataa(\Mux19~2_combout ),
	.datab(\ShiftRight0~80_combout ),
	.datac(\Mux18~4_combout ),
	.datad(\Mux18~3_combout ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hCA0F;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N18
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (\Mux18~2_combout  & (((\Mux19~3_combout )))) # (!\Mux18~2_combout  & ((\Mux19~3_combout  & (\ShiftRight0~66_combout )) # (!\Mux19~3_combout  & ((\ShiftRight0~72_combout )))))

	.dataa(\ShiftRight0~66_combout ),
	.datab(\Mux18~2_combout ),
	.datac(\Mux19~3_combout ),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hE3E0;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N30
cycloneive_lcell_comb \ShiftRight0~81 (
// Equation(s):
// \ShiftRight0~81_combout  = (!\Mux2~2_combout  & \ShiftRight0~61_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux2~2_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~81 .lut_mask = 16'h0F00;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N20
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (\Mux18~4_combout  & (((\ShiftRight0~81_combout  & \Mux18~3_combout )))) # (!\Mux18~4_combout  & ((\Mux18~5_combout ) # ((!\Mux18~3_combout ))))

	.dataa(\Mux18~5_combout ),
	.datab(\ShiftRight0~81_combout ),
	.datac(\Mux18~4_combout ),
	.datad(\Mux18~3_combout ),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hCA0F;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N2
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (\Mux18~2_combout  & (((\Mux18~6_combout )))) # (!\Mux18~2_combout  & ((\Mux18~6_combout  & ((\ShiftRight0~49_combout ))) # (!\Mux18~6_combout  & (\ShiftRight0~59_combout ))))

	.dataa(\Mux18~2_combout ),
	.datab(\ShiftRight0~59_combout ),
	.datac(\ShiftRight0~49_combout ),
	.datad(\Mux18~6_combout ),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hFA44;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N18
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (\Mux0~4_combout  & ((\Selector97~2_combout  & ((\ShiftLeft0~24_combout ))) # (!\Selector97~2_combout  & (\ShiftLeft0~31_combout ))))

	.dataa(Selector971),
	.datab(\Mux0~4_combout ),
	.datac(\ShiftLeft0~31_combout ),
	.datad(\ShiftLeft0~24_combout ),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hC840;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N0
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (\Mux18~3_combout  & ((\Mux18~4_combout  & (\ShiftRight0~103_combout )) # (!\Mux18~4_combout  & ((\Mux17~2_combout ))))) # (!\Mux18~3_combout  & (((!\Mux18~4_combout ))))

	.dataa(\ShiftRight0~103_combout ),
	.datab(\Mux18~3_combout ),
	.datac(\Mux18~4_combout ),
	.datad(\Mux17~2_combout ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'h8F83;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N10
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (\Mux18~2_combout  & (((\Mux17~3_combout )))) # (!\Mux18~2_combout  & ((\Mux17~3_combout  & ((\ShiftRight0~36_combout ))) # (!\Mux17~3_combout  & (\ShiftRight0~43_combout ))))

	.dataa(\ShiftRight0~43_combout ),
	.datab(\ShiftRight0~36_combout ),
	.datac(\Mux18~2_combout ),
	.datad(\Mux17~3_combout ),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hFC0A;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N10
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (\Mux0~4_combout  & ((\Selector97~2_combout  & (\ShiftLeft0~47_combout )) # (!\Selector97~2_combout  & ((\ShiftLeft0~52_combout )))))

	.dataa(Selector971),
	.datab(\Mux0~4_combout ),
	.datac(\ShiftLeft0~47_combout ),
	.datad(\ShiftLeft0~52_combout ),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hC480;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N28
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (\Mux18~4_combout  & (\Mux18~3_combout  & (\ShiftRight0~7_combout ))) # (!\Mux18~4_combout  & (((\Mux16~2_combout )) # (!\Mux18~3_combout )))

	.dataa(\Mux18~4_combout ),
	.datab(\Mux18~3_combout ),
	.datac(\ShiftRight0~7_combout ),
	.datad(\Mux16~2_combout ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hD591;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N6
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (\Mux18~2_combout  & (((\Mux16~3_combout )))) # (!\Mux18~2_combout  & ((\Mux16~3_combout  & (\ShiftRight0~14_combout )) # (!\Mux16~3_combout  & ((\ShiftRight0~28_combout )))))

	.dataa(\ShiftRight0~14_combout ),
	.datab(\Mux18~2_combout ),
	.datac(\ShiftRight0~28_combout ),
	.datad(\Mux16~3_combout ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hEE30;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N14
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (\Selector98~2_combout  & (Selector2 $ (((Selector3) # (Mux29))))) # (!\Selector98~2_combout  & ((Selector2 & (Selector3 $ (Mux29))) # (!Selector2 & (Selector3 & Mux29))))

	.dataa(Selector2),
	.datab(Selector981),
	.datac(Selector3),
	.datad(Mux29),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'h5668;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N26
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (Selector3 & !Selector2)

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector3),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'h00F0;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N0
cycloneive_lcell_comb \ShiftRight0~91 (
// Equation(s):
// \ShiftRight0~91_combout  = (\Selector97~2_combout  & (\ShiftRight0~77_combout )) # (!\Selector97~2_combout  & ((\ShiftRight0~86_combout )))

	.dataa(Selector971),
	.datab(gnd),
	.datac(\ShiftRight0~77_combout ),
	.datad(\ShiftRight0~86_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~91 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N20
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (Selector2) # ((Selector3 & \Selector96~2_combout ))

	.dataa(gnd),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector961),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hFCCC;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N20
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (Selector2) # ((!Selector3 & \Mux0~4_combout ))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\Mux0~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hBABA;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N18
cycloneive_lcell_comb \ShiftLeft0~92 (
// Equation(s):
// \ShiftLeft0~92_combout  = (!\Mux2~2_combout  & \ShiftLeft0~20_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux2~2_combout ),
	.datad(\ShiftLeft0~20_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~92 .lut_mask = 16'h0F00;
defparam \ShiftLeft0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N22
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (\Mux28~1_combout  & ((\Add0~37_combout ) # ((!\Mux28~0_combout )))) # (!\Mux28~1_combout  & (((\Mux28~0_combout  & \ShiftLeft0~92_combout ))))

	.dataa(\Add0~37_combout ),
	.datab(\Mux28~1_combout ),
	.datac(\Mux28~0_combout ),
	.datad(\ShiftLeft0~92_combout ),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hBC8C;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N26
cycloneive_lcell_comb \ShiftRight0~68 (
// Equation(s):
// \ShiftRight0~68_combout  = (\Selector100~4_combout  & ((Mux26))) # (!\Selector100~4_combout  & (Mux27))

	.dataa(gnd),
	.datab(Mux27),
	.datac(Mux26),
	.datad(Selector1002),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~68 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N30
cycloneive_lcell_comb \ShiftRight0~90 (
// Equation(s):
// \ShiftRight0~90_combout  = (\Selector100~4_combout  & ((Mux28))) # (!\Selector100~4_combout  & (Mux29))

	.dataa(Selector1002),
	.datab(Mux29),
	.datac(gnd),
	.datad(Mux28),
	.cin(gnd),
	.combout(\ShiftRight0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~90 .lut_mask = 16'hEE44;
defparam \ShiftRight0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N10
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (\Mux2~2_combout  & ((\ShiftRight0~38_combout ) # ((\Mux2~1_combout )))) # (!\Mux2~2_combout  & (((\ShiftRight0~90_combout  & !\Mux2~1_combout ))))

	.dataa(\ShiftRight0~38_combout ),
	.datab(\Mux2~2_combout ),
	.datac(\ShiftRight0~90_combout ),
	.datad(\Mux2~1_combout ),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hCCB8;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N12
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (\Mux2~1_combout  & ((\Mux29~0_combout  & ((\ShiftRight0~87_combout ))) # (!\Mux29~0_combout  & (\ShiftRight0~68_combout )))) # (!\Mux2~1_combout  & (((\Mux29~0_combout ))))

	.dataa(\Mux2~1_combout ),
	.datab(\ShiftRight0~68_combout ),
	.datac(\ShiftRight0~87_combout ),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hF588;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N8
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (\Mux6~17_combout  & ((\Mux29~2_combout  & (\ShiftRight0~91_combout )) # (!\Mux29~2_combout  & ((\Mux29~1_combout ))))) # (!\Mux6~17_combout  & (((\Mux29~2_combout ))))

	.dataa(\Mux6~17_combout ),
	.datab(\ShiftRight0~91_combout ),
	.datac(\Mux29~2_combout ),
	.datad(\Mux29~1_combout ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hDAD0;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N0
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (!Selector0 & (!Selector1 & ((!\ShiftLeft0~32_combout ) # (!\Mux6~17_combout ))))

	.dataa(Selector0),
	.datab(Selector1),
	.datac(\Mux6~17_combout ),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'h0111;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N16
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (\Selector97~2_combout  & (Selector2 $ (((Selector3) # (Mux28))))) # (!\Selector97~2_combout  & ((Selector2 & (Selector3 $ (Mux28))) # (!Selector2 & (Selector3 & Mux28))))

	.dataa(Selector971),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Mux28),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'h3668;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N30
cycloneive_lcell_comb \ShiftRight0~92 (
// Equation(s):
// \ShiftRight0~92_combout  = (\Selector100~4_combout  & (Mux27)) # (!\Selector100~4_combout  & ((Mux28)))

	.dataa(gnd),
	.datab(Mux27),
	.datac(Mux28),
	.datad(Selector1002),
	.cin(gnd),
	.combout(\ShiftRight0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~92 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N28
cycloneive_lcell_comb \ShiftRight0~19 (
// Equation(s):
// \ShiftRight0~19_combout  = (\Selector99~2_combout  & ((Mux22))) # (!\Selector99~2_combout  & (Mux24))

	.dataa(Mux24),
	.datab(Selector991),
	.datac(gnd),
	.datad(Mux22),
	.cin(gnd),
	.combout(\ShiftRight0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~19 .lut_mask = 16'hEE22;
defparam \ShiftRight0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N2
cycloneive_lcell_comb \ShiftRight0~20 (
// Equation(s):
// \ShiftRight0~20_combout  = (\Selector100~4_combout  & (\ShiftRight0~18_combout )) # (!\Selector100~4_combout  & ((\ShiftRight0~19_combout )))

	.dataa(Selector1002),
	.datab(gnd),
	.datac(\ShiftRight0~18_combout ),
	.datad(\ShiftRight0~19_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~20 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N30
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (\Mux2~1_combout  & (\Mux2~2_combout )) # (!\Mux2~1_combout  & ((\Mux2~2_combout  & ((\ShiftRight0~20_combout ))) # (!\Mux2~2_combout  & (\ShiftRight0~92_combout ))))

	.dataa(\Mux2~1_combout ),
	.datab(\Mux2~2_combout ),
	.datac(\ShiftRight0~92_combout ),
	.datad(\ShiftRight0~20_combout ),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hDC98;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N6
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (\Mux2~1_combout  & ((\Mux28~2_combout  & ((\ShiftRight0~89_combout ))) # (!\Mux28~2_combout  & (\ShiftRight0~53_combout )))) # (!\Mux2~1_combout  & (((\Mux28~2_combout ))))

	.dataa(\ShiftRight0~53_combout ),
	.datab(\Mux2~1_combout ),
	.datac(\Mux28~2_combout ),
	.datad(\ShiftRight0~89_combout ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hF838;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N18
cycloneive_lcell_comb \ShiftLeft0~93 (
// Equation(s):
// \ShiftLeft0~93_combout  = (!\Mux2~2_combout  & ((\ShiftLeft0~42_combout ) # ((\Selector99~2_combout  & \ShiftLeft0~43_combout ))))

	.dataa(\ShiftLeft0~42_combout ),
	.datab(\Mux2~2_combout ),
	.datac(Selector991),
	.datad(\ShiftLeft0~43_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~93 .lut_mask = 16'h3222;
defparam \ShiftLeft0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N4
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (\Mux28~1_combout  & ((\Add0~39_combout ) # ((!\Mux28~0_combout )))) # (!\Mux28~1_combout  & (((\Mux28~0_combout  & \ShiftLeft0~93_combout ))))

	.dataa(\Add0~39_combout ),
	.datab(\Mux28~1_combout ),
	.datac(\Mux28~0_combout ),
	.datad(\ShiftLeft0~93_combout ),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hBC8C;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N26
cycloneive_lcell_comb \ShiftRight0~93 (
// Equation(s):
// \ShiftRight0~93_combout  = (\Selector97~2_combout  & ((\ShiftRight0~76_combout ))) # (!\Selector97~2_combout  & (\ShiftRight0~88_combout ))

	.dataa(gnd),
	.datab(Selector971),
	.datac(\ShiftRight0~88_combout ),
	.datad(\ShiftRight0~76_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~93 .lut_mask = 16'hFC30;
defparam \ShiftRight0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N10
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (\Mux6~17_combout  & ((\Mux28~4_combout  & ((\ShiftRight0~93_combout ))) # (!\Mux28~4_combout  & (\Mux28~3_combout )))) # (!\Mux6~17_combout  & (((\Mux28~4_combout ))))

	.dataa(\Mux28~3_combout ),
	.datab(\Mux6~17_combout ),
	.datac(\Mux28~4_combout ),
	.datad(\ShiftRight0~93_combout ),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hF838;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N18
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (Selector3 & (Selector2 $ (((\Selector77~1_combout ) # (Mux8))))) # (!Selector3 & ((Selector2 & (\Selector77~1_combout  $ (Mux8))) # (!Selector2 & (\Selector77~1_combout  & Mux8))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(Selector771),
	.datad(Mux8),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'h5668;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N12
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (!Selector0 & (Selector1 & \Mux8~4_combout ))

	.dataa(gnd),
	.datab(Selector0),
	.datac(Selector1),
	.datad(\Mux8~4_combout ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'h3000;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N0
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (Selector3) # ((\Selector97~2_combout  & \Mux0~4_combout ))

	.dataa(gnd),
	.datab(Selector971),
	.datac(Selector3),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hFCF0;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N14
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (\Mux0~6_combout  & ((\Mux0~7_combout  & ((\ShiftRight0~29_combout ))) # (!\Mux0~7_combout  & (\Mux8~10_combout )))) # (!\Mux0~6_combout  & (((!\Mux0~7_combout ))))

	.dataa(\Mux8~10_combout ),
	.datab(\Mux0~6_combout ),
	.datac(\ShiftRight0~29_combout ),
	.datad(\Mux0~7_combout ),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hC0BB;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N8
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (\Mux0~5_combout  & (((\Mux8~6_combout )))) # (!\Mux0~5_combout  & ((\Mux8~6_combout  & (\ShiftLeft0~37_combout )) # (!\Mux8~6_combout  & ((\ShiftLeft0~52_combout )))))

	.dataa(\ShiftLeft0~37_combout ),
	.datab(\Mux0~5_combout ),
	.datac(\Mux8~6_combout ),
	.datad(\ShiftLeft0~52_combout ),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hE3E0;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N16
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// \Mux8~9_combout  = (Selector2 & (!Selector0 & (!Selector1 & \Add0~79_combout )))

	.dataa(Selector2),
	.datab(Selector0),
	.datac(Selector1),
	.datad(\Add0~79_combout ),
	.cin(gnd),
	.combout(\Mux8~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'h0200;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N14
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (!\Selector97~2_combout  & (!\ShiftLeft0~18_combout  & (!\ShiftLeft0~16_combout  & !\ShiftLeft0~15_combout )))

	.dataa(Selector971),
	.datab(\ShiftLeft0~18_combout ),
	.datac(\ShiftLeft0~16_combout ),
	.datad(\ShiftLeft0~15_combout ),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'h0001;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N30
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (\Mux15~2_combout  & \ShiftLeft0~55_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux15~2_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hF000;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N20
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (\Mux0~6_combout  & ((\Mux0~7_combout  & (\ShiftRight0~62_combout )) # (!\Mux0~7_combout  & ((\Mux10~2_combout ))))) # (!\Mux0~6_combout  & (((!\Mux0~7_combout ))))

	.dataa(\ShiftRight0~62_combout ),
	.datab(\Mux0~6_combout ),
	.datac(\Mux10~2_combout ),
	.datad(\Mux0~7_combout ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'h88F3;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N26
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (\Mux0~5_combout  & (((\Mux10~3_combout )))) # (!\Mux0~5_combout  & ((\Mux10~3_combout  & ((\ShiftLeft0~91_combout ))) # (!\Mux10~3_combout  & (\ShiftLeft0~90_combout ))))

	.dataa(\ShiftLeft0~90_combout ),
	.datab(\ShiftLeft0~91_combout ),
	.datac(\Mux0~5_combout ),
	.datad(\Mux10~3_combout ),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hFC0A;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N0
cycloneive_lcell_comb \Add0~9 (
// Equation(s):
// \Add0~9_combout  = Selector3 $ (((\Selector79~0_combout ) # ((\Selector95~0_combout  & Mux42))))

	.dataa(Selector95),
	.datab(Mux42),
	.datac(Selector3),
	.datad(Selector79),
	.cin(gnd),
	.combout(\Add0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~9 .lut_mask = 16'h0F78;
defparam \Add0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N6
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = Selector3 $ (((\Selector78~0_combout ) # ((\Selector95~0_combout  & Mux41))))

	.dataa(Selector95),
	.datab(Selector3),
	.datac(Selector78),
	.datad(Mux41),
	.cin(gnd),
	.combout(\Add0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h363C;
defparam \Add0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N10
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (\Mux0~6_combout  & ((\Mux0~7_combout  & ((\ShiftRight0~44_combout ))) # (!\Mux0~7_combout  & (\Mux9~8_combout )))) # (!\Mux0~6_combout  & (((!\Mux0~7_combout ))))

	.dataa(\Mux9~8_combout ),
	.datab(\Mux0~6_combout ),
	.datac(\ShiftRight0~44_combout ),
	.datad(\Mux0~7_combout ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hC0BB;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N20
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (\Mux0~5_combout  & (((\Mux9~4_combout )))) # (!\Mux0~5_combout  & ((\Mux9~4_combout  & ((\ShiftLeft0~6_combout ))) # (!\Mux9~4_combout  & (\ShiftLeft0~31_combout ))))

	.dataa(\Mux0~5_combout ),
	.datab(\ShiftLeft0~31_combout ),
	.datac(\ShiftLeft0~6_combout ),
	.datad(\Mux9~4_combout ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hFA44;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N8
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (\Selector99~2_combout  & (Selector2 $ (((Mux30) # (Selector3))))) # (!\Selector99~2_combout  & ((Selector2 & (Mux30 $ (Selector3))) # (!Selector2 & (Mux30 & Selector3))))

	.dataa(Selector991),
	.datab(Selector2),
	.datac(Mux30),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'h3668;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N10
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (Selector1 & (((\Mux30~3_combout )))) # (!Selector1 & (Selector2 & ((\Add0~35_combout ))))

	.dataa(Selector2),
	.datab(Selector1),
	.datac(\Mux30~3_combout ),
	.datad(\Add0~35_combout ),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hE2C0;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N8
cycloneive_lcell_comb \ShiftRight0~94 (
// Equation(s):
// \ShiftRight0~94_combout  = (!\Selector99~2_combout  & ((\Selector100~4_combout  & ((Mux29))) # (!\Selector100~4_combout  & (Mux30))))

	.dataa(Selector1002),
	.datab(Selector991),
	.datac(Mux30),
	.datad(Mux29),
	.cin(gnd),
	.combout(\ShiftRight0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~94 .lut_mask = 16'h3210;
defparam \ShiftRight0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N30
cycloneive_lcell_comb \ShiftRight0~95 (
// Equation(s):
// \ShiftRight0~95_combout  = (!\Selector98~2_combout  & ((\ShiftRight0~94_combout ) # ((\Selector99~2_combout  & \ShiftRight0~92_combout ))))

	.dataa(Selector991),
	.datab(\ShiftRight0~94_combout ),
	.datac(Selector981),
	.datad(\ShiftRight0~92_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~95 .lut_mask = 16'h0E0C;
defparam \ShiftRight0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N12
cycloneive_lcell_comb \ShiftRight0~96 (
// Equation(s):
// \ShiftRight0~96_combout  = (!\Selector97~2_combout  & ((\ShiftRight0~95_combout ) # ((\Selector98~2_combout  & \ShiftRight0~54_combout ))))

	.dataa(Selector981),
	.datab(Selector971),
	.datac(\ShiftRight0~95_combout ),
	.datad(\ShiftRight0~54_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~96 .lut_mask = 16'h3230;
defparam \ShiftRight0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N26
cycloneive_lcell_comb \ShiftRight0~97 (
// Equation(s):
// \ShiftRight0~97_combout  = (!\Selector96~2_combout  & ((\ShiftRight0~96_combout ) # ((\Selector97~2_combout  & \ShiftRight0~85_combout ))))

	.dataa(Selector971),
	.datab(Selector961),
	.datac(\ShiftRight0~85_combout ),
	.datad(\ShiftRight0~96_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~97 .lut_mask = 16'h3320;
defparam \ShiftRight0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N16
cycloneive_lcell_comb \ShiftRight0~98 (
// Equation(s):
// \ShiftRight0~98_combout  = (\Selector98~2_combout  & (\ShiftRight0~61_combout )) # (!\Selector98~2_combout  & ((\ShiftRight0~56_combout )))

	.dataa(\ShiftRight0~61_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~56_combout ),
	.datad(Selector981),
	.cin(gnd),
	.combout(\ShiftRight0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~98 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N18
cycloneive_lcell_comb \ShiftRight0~99 (
// Equation(s):
// \ShiftRight0~99_combout  = (\Selector97~2_combout  & ((\ShiftRight0~98_combout ))) # (!\Selector97~2_combout  & (\ShiftRight0~84_combout ))

	.dataa(\ShiftRight0~84_combout ),
	.datab(gnd),
	.datac(Selector971),
	.datad(\ShiftRight0~98_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~99 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N0
cycloneive_lcell_comb \ShiftRight0~100 (
// Equation(s):
// \ShiftRight0~100_combout  = (\ShiftRight0~97_combout ) # ((\Selector96~2_combout  & \ShiftRight0~99_combout ))

	.dataa(gnd),
	.datab(Selector961),
	.datac(\ShiftRight0~97_combout ),
	.datad(\ShiftRight0~99_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~100 .lut_mask = 16'hFCF0;
defparam \ShiftRight0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N22
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (Selector3 & (!\ShiftLeft0~32_combout  & (\Mux30~0_combout  & \ShiftRight0~100_combout )))

	.dataa(Selector3),
	.datab(\ShiftLeft0~32_combout ),
	.datac(\Mux30~0_combout ),
	.datad(\ShiftRight0~100_combout ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'h2000;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N14
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (!\Selector98~2_combout  & (!\Selector99~2_combout  & (\ShiftLeft0~43_combout  & \Mux15~2_combout )))

	.dataa(Selector981),
	.datab(Selector991),
	.datac(\ShiftLeft0~43_combout ),
	.datad(\Mux15~2_combout ),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'h1000;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N28
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (\Mux30~0_combout  & (!\Selector96~2_combout  & (\Mux14~8_combout  & !Selector3)))

	.dataa(\Mux30~0_combout ),
	.datab(Selector961),
	.datac(\Mux14~8_combout ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'h0020;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N8
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = Selector3 $ (((\Selector84~1_combout ) # ((Mux47 & \Selector95~0_combout ))))

	.dataa(Mux47),
	.datab(Selector3),
	.datac(Selector84),
	.datad(Selector95),
	.cin(gnd),
	.combout(\Add0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h363C;
defparam \Add0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N4
cycloneive_lcell_comb \ShiftRight0~101 (
// Equation(s):
// \ShiftRight0~101_combout  = (\Selector98~2_combout  & ((\ShiftRight0~74_combout ))) # (!\Selector98~2_combout  & (\ShiftRight0~70_combout ))

	.dataa(gnd),
	.datab(Selector981),
	.datac(\ShiftRight0~70_combout ),
	.datad(\ShiftRight0~74_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~101 .lut_mask = 16'hFC30;
defparam \ShiftRight0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N10
cycloneive_lcell_comb \ShiftRight0~102 (
// Equation(s):
// \ShiftRight0~102_combout  = (\Selector97~2_combout  & (\ShiftRight0~101_combout )) # (!\Selector97~2_combout  & ((\ShiftRight0~82_combout )))

	.dataa(gnd),
	.datab(Selector971),
	.datac(\ShiftRight0~101_combout ),
	.datad(\ShiftRight0~82_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~102 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N28
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (\Mux0~6_combout  & ((\Mux0~7_combout  & ((\ShiftRight0~102_combout ))) # (!\Mux0~7_combout  & (\Mux15~3_combout )))) # (!\Mux0~6_combout  & (((!\Mux0~7_combout ))))

	.dataa(\Mux15~3_combout ),
	.datab(\Mux0~6_combout ),
	.datac(\Mux0~7_combout ),
	.datad(\ShiftRight0~102_combout ),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hCB0B;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N18
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (\Mux0~5_combout  & (((\Mux15~4_combout )))) # (!\Mux0~5_combout  & ((\Mux15~4_combout  & (\ShiftLeft0~83_combout )) # (!\Mux15~4_combout  & ((\ShiftLeft0~86_combout )))))

	.dataa(\ShiftLeft0~83_combout ),
	.datab(\ShiftLeft0~86_combout ),
	.datac(\Mux0~5_combout ),
	.datad(\Mux15~4_combout ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hFA0C;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N24
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (\Mux0~6_combout  & ((\Mux0~7_combout  & ((\ShiftRight0~99_combout ))) # (!\Mux0~7_combout  & (\Mux14~8_combout )))) # (!\Mux0~6_combout  & (!\Mux0~7_combout ))

	.dataa(\Mux0~6_combout ),
	.datab(\Mux0~7_combout ),
	.datac(\Mux14~8_combout ),
	.datad(\ShiftRight0~99_combout ),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hB931;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N18
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (\Mux0~5_combout  & (((\Mux14~4_combout )))) # (!\Mux0~5_combout  & ((\Mux14~4_combout  & ((\ShiftLeft0~70_combout ))) # (!\Mux14~4_combout  & (\ShiftLeft0~78_combout ))))

	.dataa(\ShiftLeft0~78_combout ),
	.datab(\Mux0~5_combout ),
	.datac(\ShiftLeft0~70_combout ),
	.datad(\Mux14~4_combout ),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hFC22;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N12
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = Selector3 $ (((\Selector82~0_combout ) # ((Mux45 & \Selector95~0_combout ))))

	.dataa(Mux45),
	.datab(Selector95),
	.datac(Selector3),
	.datad(Selector82),
	.cin(gnd),
	.combout(\Add0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h0F78;
defparam \Add0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N2
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (\ShiftLeft0~20_combout  & (!\Mux2~2_combout  & !\ShiftLeft0~32_combout ))

	.dataa(\ShiftLeft0~20_combout ),
	.datab(gnd),
	.datac(\Mux2~2_combout ),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'h000A;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N24
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (\Mux0~6_combout  & ((\Mux0~7_combout  & (\ShiftRight0~91_combout )) # (!\Mux0~7_combout  & ((\Mux13~2_combout ))))) # (!\Mux0~6_combout  & (((!\Mux0~7_combout ))))

	.dataa(\Mux0~6_combout ),
	.datab(\ShiftRight0~91_combout ),
	.datac(\Mux13~2_combout ),
	.datad(\Mux0~7_combout ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'h88F5;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N2
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (\Mux0~5_combout  & (((\Mux13~3_combout )))) # (!\Mux0~5_combout  & ((\Mux13~3_combout  & ((\ShiftLeft0~63_combout ))) # (!\Mux13~3_combout  & (\ShiftLeft0~64_combout ))))

	.dataa(\ShiftLeft0~64_combout ),
	.datab(\Mux0~5_combout ),
	.datac(\ShiftLeft0~63_combout ),
	.datad(\Mux13~3_combout ),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hFC22;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N22
cycloneive_lcell_comb \Add0~11 (
// Equation(s):
// \Add0~11_combout  = Selector3 $ (((\Selector81~0_combout ) # ((\Selector95~0_combout  & Mux44))))

	.dataa(Selector95),
	.datab(Selector81),
	.datac(Selector3),
	.datad(Mux44),
	.cin(gnd),
	.combout(\Add0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~11 .lut_mask = 16'h1E3C;
defparam \Add0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N8
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (!\Mux2~2_combout  & (\ShiftLeft0~44_combout  & !\ShiftLeft0~32_combout ))

	.dataa(\Mux2~2_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~44_combout ),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'h0050;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N10
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (\Mux0~6_combout  & ((\Mux0~7_combout  & (\ShiftRight0~93_combout )) # (!\Mux0~7_combout  & ((\Mux12~2_combout ))))) # (!\Mux0~6_combout  & (((!\Mux0~7_combout ))))

	.dataa(\ShiftRight0~93_combout ),
	.datab(\Mux0~6_combout ),
	.datac(\Mux12~2_combout ),
	.datad(\Mux0~7_combout ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'h88F3;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N28
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (\Mux0~5_combout  & (((\Mux12~3_combout )))) # (!\Mux0~5_combout  & ((\Mux12~3_combout  & ((\ShiftLeft0~60_combout ))) # (!\Mux12~3_combout  & (\ShiftLeft0~61_combout ))))

	.dataa(\ShiftLeft0~61_combout ),
	.datab(\Mux0~5_combout ),
	.datac(\ShiftLeft0~60_combout ),
	.datad(\Mux12~3_combout ),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hFC22;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N18
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = Selector3 $ (((\Selector80~0_combout ) # ((Mux43 & \Selector95~0_combout ))))

	.dataa(Mux43),
	.datab(Selector3),
	.datac(Selector80),
	.datad(Selector95),
	.cin(gnd),
	.combout(\Add0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h363C;
defparam \Add0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N0
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (\Mux0~6_combout  & ((\Mux0~7_combout  & ((\ShiftRight0~75_combout ))) # (!\Mux0~7_combout  & (\Mux11~2_combout )))) # (!\Mux0~6_combout  & (((!\Mux0~7_combout ))))

	.dataa(\Mux11~2_combout ),
	.datab(\Mux0~6_combout ),
	.datac(\ShiftRight0~75_combout ),
	.datad(\Mux0~7_combout ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hC0BB;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N2
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (\Mux0~5_combout  & (((\Mux11~3_combout )))) # (!\Mux0~5_combout  & ((\Mux11~3_combout  & ((\ShiftLeft0~89_combout ))) # (!\Mux11~3_combout  & (\ShiftLeft0~88_combout ))))

	.dataa(\ShiftLeft0~88_combout ),
	.datab(\ShiftLeft0~89_combout ),
	.datac(\Mux0~5_combout ),
	.datad(\Mux11~3_combout ),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hFC0A;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N30
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (Selector0 & (Selector2 & !Selector1))

	.dataa(gnd),
	.datab(Selector0),
	.datac(Selector2),
	.datad(Selector1),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'h00C0;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N0
cycloneive_lcell_comb \LessThan0~1 (
// Equation(s):
// \LessThan0~1_cout  = CARRY((\Selector100~4_combout  & !Mux31))

	.dataa(Selector1002),
	.datab(Mux31),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
// synopsys translate_off
defparam \LessThan0~1 .lut_mask = 16'h0022;
defparam \LessThan0~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N2
cycloneive_lcell_comb \LessThan0~3 (
// Equation(s):
// \LessThan0~3_cout  = CARRY((\Selector99~2_combout  & (Mux30 & !\LessThan0~1_cout )) # (!\Selector99~2_combout  & ((Mux30) # (!\LessThan0~1_cout ))))

	.dataa(Selector991),
	.datab(Mux30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
// synopsys translate_off
defparam \LessThan0~3 .lut_mask = 16'h004D;
defparam \LessThan0~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N4
cycloneive_lcell_comb \LessThan0~5 (
// Equation(s):
// \LessThan0~5_cout  = CARRY((Mux29 & (\Selector98~2_combout  & !\LessThan0~3_cout )) # (!Mux29 & ((\Selector98~2_combout ) # (!\LessThan0~3_cout ))))

	.dataa(Mux29),
	.datab(Selector981),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
// synopsys translate_off
defparam \LessThan0~5 .lut_mask = 16'h004D;
defparam \LessThan0~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N6
cycloneive_lcell_comb \LessThan0~7 (
// Equation(s):
// \LessThan0~7_cout  = CARRY((\Selector97~2_combout  & (Mux28 & !\LessThan0~5_cout )) # (!\Selector97~2_combout  & ((Mux28) # (!\LessThan0~5_cout ))))

	.dataa(Selector971),
	.datab(Mux28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
// synopsys translate_off
defparam \LessThan0~7 .lut_mask = 16'h004D;
defparam \LessThan0~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N8
cycloneive_lcell_comb \LessThan0~9 (
// Equation(s):
// \LessThan0~9_cout  = CARRY((\Selector96~2_combout  & ((!\LessThan0~7_cout ) # (!Mux27))) # (!\Selector96~2_combout  & (!Mux27 & !\LessThan0~7_cout )))

	.dataa(Selector961),
	.datab(Mux27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
// synopsys translate_off
defparam \LessThan0~9 .lut_mask = 16'h002B;
defparam \LessThan0~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N10
cycloneive_lcell_comb \LessThan0~11 (
// Equation(s):
// \LessThan0~11_cout  = CARRY((\Selector95~3_combout  & (Mux26 & !\LessThan0~9_cout )) # (!\Selector95~3_combout  & ((Mux26) # (!\LessThan0~9_cout ))))

	.dataa(Selector952),
	.datab(Mux26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
// synopsys translate_off
defparam \LessThan0~11 .lut_mask = 16'h004D;
defparam \LessThan0~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N12
cycloneive_lcell_comb \LessThan0~13 (
// Equation(s):
// \LessThan0~13_cout  = CARRY((\Selector94~1_combout  & ((!\LessThan0~11_cout ) # (!Mux25))) # (!\Selector94~1_combout  & (!Mux25 & !\LessThan0~11_cout )))

	.dataa(Selector941),
	.datab(Mux25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
// synopsys translate_off
defparam \LessThan0~13 .lut_mask = 16'h002B;
defparam \LessThan0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N14
cycloneive_lcell_comb \LessThan0~15 (
// Equation(s):
// \LessThan0~15_cout  = CARRY((Mux24 & ((!\LessThan0~13_cout ) # (!\Selector93~1_combout ))) # (!Mux24 & (!\Selector93~1_combout  & !\LessThan0~13_cout )))

	.dataa(Mux24),
	.datab(Selector931),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
// synopsys translate_off
defparam \LessThan0~15 .lut_mask = 16'h002B;
defparam \LessThan0~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N16
cycloneive_lcell_comb \LessThan0~17 (
// Equation(s):
// \LessThan0~17_cout  = CARRY((\Selector92~1_combout  & ((!\LessThan0~15_cout ) # (!Mux23))) # (!\Selector92~1_combout  & (!Mux23 & !\LessThan0~15_cout )))

	.dataa(Selector921),
	.datab(Mux23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
// synopsys translate_off
defparam \LessThan0~17 .lut_mask = 16'h002B;
defparam \LessThan0~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N18
cycloneive_lcell_comb \LessThan0~19 (
// Equation(s):
// \LessThan0~19_cout  = CARRY((Mux22 & ((!\LessThan0~17_cout ) # (!\Selector91~1_combout ))) # (!Mux22 & (!\Selector91~1_combout  & !\LessThan0~17_cout )))

	.dataa(Mux22),
	.datab(Selector911),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
// synopsys translate_off
defparam \LessThan0~19 .lut_mask = 16'h002B;
defparam \LessThan0~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N20
cycloneive_lcell_comb \LessThan0~21 (
// Equation(s):
// \LessThan0~21_cout  = CARRY((\Selector90~1_combout  & ((!\LessThan0~19_cout ) # (!Mux21))) # (!\Selector90~1_combout  & (!Mux21 & !\LessThan0~19_cout )))

	.dataa(Selector901),
	.datab(Mux21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
// synopsys translate_off
defparam \LessThan0~21 .lut_mask = 16'h002B;
defparam \LessThan0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N22
cycloneive_lcell_comb \LessThan0~23 (
// Equation(s):
// \LessThan0~23_cout  = CARRY((\Selector89~1_combout  & (Mux20 & !\LessThan0~21_cout )) # (!\Selector89~1_combout  & ((Mux20) # (!\LessThan0~21_cout ))))

	.dataa(Selector891),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
// synopsys translate_off
defparam \LessThan0~23 .lut_mask = 16'h004D;
defparam \LessThan0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N24
cycloneive_lcell_comb \LessThan0~25 (
// Equation(s):
// \LessThan0~25_cout  = CARRY((Mux19 & (\Selector88~1_combout  & !\LessThan0~23_cout )) # (!Mux19 & ((\Selector88~1_combout ) # (!\LessThan0~23_cout ))))

	.dataa(Mux19),
	.datab(Selector881),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
// synopsys translate_off
defparam \LessThan0~25 .lut_mask = 16'h004D;
defparam \LessThan0~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N26
cycloneive_lcell_comb \LessThan0~27 (
// Equation(s):
// \LessThan0~27_cout  = CARRY((\Selector87~1_combout  & (Mux18 & !\LessThan0~25_cout )) # (!\Selector87~1_combout  & ((Mux18) # (!\LessThan0~25_cout ))))

	.dataa(Selector871),
	.datab(Mux18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
// synopsys translate_off
defparam \LessThan0~27 .lut_mask = 16'h004D;
defparam \LessThan0~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N28
cycloneive_lcell_comb \LessThan0~29 (
// Equation(s):
// \LessThan0~29_cout  = CARRY((\Selector86~1_combout  & ((!\LessThan0~27_cout ) # (!Mux17))) # (!\Selector86~1_combout  & (!Mux17 & !\LessThan0~27_cout )))

	.dataa(Selector861),
	.datab(Mux17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
// synopsys translate_off
defparam \LessThan0~29 .lut_mask = 16'h002B;
defparam \LessThan0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N30
cycloneive_lcell_comb \LessThan0~31 (
// Equation(s):
// \LessThan0~31_cout  = CARRY((\Selector85~1_combout  & (Mux16 & !\LessThan0~29_cout )) # (!\Selector85~1_combout  & ((Mux16) # (!\LessThan0~29_cout ))))

	.dataa(Selector851),
	.datab(Mux16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
// synopsys translate_off
defparam \LessThan0~31 .lut_mask = 16'h004D;
defparam \LessThan0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N0
cycloneive_lcell_comb \LessThan0~33 (
// Equation(s):
// \LessThan0~33_cout  = CARRY((Mux15 & (\Selector84~2_combout  & !\LessThan0~31_cout )) # (!Mux15 & ((\Selector84~2_combout ) # (!\LessThan0~31_cout ))))

	.dataa(Mux15),
	.datab(Selector841),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
// synopsys translate_off
defparam \LessThan0~33 .lut_mask = 16'h004D;
defparam \LessThan0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N2
cycloneive_lcell_comb \LessThan0~35 (
// Equation(s):
// \LessThan0~35_cout  = CARRY((\Selector83~1_combout  & (Mux14 & !\LessThan0~33_cout )) # (!\Selector83~1_combout  & ((Mux14) # (!\LessThan0~33_cout ))))

	.dataa(Selector831),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~33_cout ),
	.combout(),
	.cout(\LessThan0~35_cout ));
// synopsys translate_off
defparam \LessThan0~35 .lut_mask = 16'h004D;
defparam \LessThan0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N4
cycloneive_lcell_comb \LessThan0~37 (
// Equation(s):
// \LessThan0~37_cout  = CARRY((Mux13 & (\Selector82~1_combout  & !\LessThan0~35_cout )) # (!Mux13 & ((\Selector82~1_combout ) # (!\LessThan0~35_cout ))))

	.dataa(Mux13),
	.datab(Selector821),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~35_cout ),
	.combout(),
	.cout(\LessThan0~37_cout ));
// synopsys translate_off
defparam \LessThan0~37 .lut_mask = 16'h004D;
defparam \LessThan0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N6
cycloneive_lcell_comb \LessThan0~39 (
// Equation(s):
// \LessThan0~39_cout  = CARRY((Mux12 & ((!\LessThan0~37_cout ) # (!\Selector81~1_combout ))) # (!Mux12 & (!\Selector81~1_combout  & !\LessThan0~37_cout )))

	.dataa(Mux12),
	.datab(Selector811),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~37_cout ),
	.combout(),
	.cout(\LessThan0~39_cout ));
// synopsys translate_off
defparam \LessThan0~39 .lut_mask = 16'h002B;
defparam \LessThan0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N8
cycloneive_lcell_comb \LessThan0~41 (
// Equation(s):
// \LessThan0~41_cout  = CARRY((\Selector80~1_combout  & ((!\LessThan0~39_cout ) # (!Mux11))) # (!\Selector80~1_combout  & (!Mux11 & !\LessThan0~39_cout )))

	.dataa(Selector801),
	.datab(Mux11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~39_cout ),
	.combout(),
	.cout(\LessThan0~41_cout ));
// synopsys translate_off
defparam \LessThan0~41 .lut_mask = 16'h002B;
defparam \LessThan0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N10
cycloneive_lcell_comb \LessThan0~43 (
// Equation(s):
// \LessThan0~43_cout  = CARRY((Mux10 & ((!\LessThan0~41_cout ) # (!\Selector79~1_combout ))) # (!Mux10 & (!\Selector79~1_combout  & !\LessThan0~41_cout )))

	.dataa(Mux10),
	.datab(Selector791),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~41_cout ),
	.combout(),
	.cout(\LessThan0~43_cout ));
// synopsys translate_off
defparam \LessThan0~43 .lut_mask = 16'h002B;
defparam \LessThan0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N12
cycloneive_lcell_comb \LessThan0~45 (
// Equation(s):
// \LessThan0~45_cout  = CARRY((\Selector78~1_combout  & ((!\LessThan0~43_cout ) # (!Mux9))) # (!\Selector78~1_combout  & (!Mux9 & !\LessThan0~43_cout )))

	.dataa(Selector781),
	.datab(Mux9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~43_cout ),
	.combout(),
	.cout(\LessThan0~45_cout ));
// synopsys translate_off
defparam \LessThan0~45 .lut_mask = 16'h002B;
defparam \LessThan0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N14
cycloneive_lcell_comb \LessThan0~47 (
// Equation(s):
// \LessThan0~47_cout  = CARRY((Mux8 & ((!\LessThan0~45_cout ) # (!\Selector77~1_combout ))) # (!Mux8 & (!\Selector77~1_combout  & !\LessThan0~45_cout )))

	.dataa(Mux8),
	.datab(Selector771),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~45_cout ),
	.combout(),
	.cout(\LessThan0~47_cout ));
// synopsys translate_off
defparam \LessThan0~47 .lut_mask = 16'h002B;
defparam \LessThan0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N16
cycloneive_lcell_comb \LessThan0~49 (
// Equation(s):
// \LessThan0~49_cout  = CARRY((Mux7 & (\Selector76~1_combout  & !\LessThan0~47_cout )) # (!Mux7 & ((\Selector76~1_combout ) # (!\LessThan0~47_cout ))))

	.dataa(Mux7),
	.datab(Selector761),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~47_cout ),
	.combout(),
	.cout(\LessThan0~49_cout ));
// synopsys translate_off
defparam \LessThan0~49 .lut_mask = 16'h004D;
defparam \LessThan0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N18
cycloneive_lcell_comb \LessThan0~51 (
// Equation(s):
// \LessThan0~51_cout  = CARRY((Mux6 & ((!\LessThan0~49_cout ) # (!\Selector75~1_combout ))) # (!Mux6 & (!\Selector75~1_combout  & !\LessThan0~49_cout )))

	.dataa(Mux6),
	.datab(Selector751),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~49_cout ),
	.combout(),
	.cout(\LessThan0~51_cout ));
// synopsys translate_off
defparam \LessThan0~51 .lut_mask = 16'h002B;
defparam \LessThan0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N20
cycloneive_lcell_comb \LessThan0~53 (
// Equation(s):
// \LessThan0~53_cout  = CARRY((\Selector74~1_combout  & ((!\LessThan0~51_cout ) # (!Mux5))) # (!\Selector74~1_combout  & (!Mux5 & !\LessThan0~51_cout )))

	.dataa(Selector741),
	.datab(Mux5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~51_cout ),
	.combout(),
	.cout(\LessThan0~53_cout ));
// synopsys translate_off
defparam \LessThan0~53 .lut_mask = 16'h002B;
defparam \LessThan0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N22
cycloneive_lcell_comb \LessThan0~55 (
// Equation(s):
// \LessThan0~55_cout  = CARRY((\Selector73~1_combout  & (Mux4 & !\LessThan0~53_cout )) # (!\Selector73~1_combout  & ((Mux4) # (!\LessThan0~53_cout ))))

	.dataa(Selector731),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~53_cout ),
	.combout(),
	.cout(\LessThan0~55_cout ));
// synopsys translate_off
defparam \LessThan0~55 .lut_mask = 16'h004D;
defparam \LessThan0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N24
cycloneive_lcell_comb \LessThan0~57 (
// Equation(s):
// \LessThan0~57_cout  = CARRY((\Selector72~1_combout  & ((!\LessThan0~55_cout ) # (!Mux3))) # (!\Selector72~1_combout  & (!Mux3 & !\LessThan0~55_cout )))

	.dataa(Selector721),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~55_cout ),
	.combout(),
	.cout(\LessThan0~57_cout ));
// synopsys translate_off
defparam \LessThan0~57 .lut_mask = 16'h002B;
defparam \LessThan0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N26
cycloneive_lcell_comb \LessThan0~59 (
// Equation(s):
// \LessThan0~59_cout  = CARRY((\Selector71~1_combout  & (Mux2 & !\LessThan0~57_cout )) # (!\Selector71~1_combout  & ((Mux2) # (!\LessThan0~57_cout ))))

	.dataa(Selector711),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~57_cout ),
	.combout(),
	.cout(\LessThan0~59_cout ));
// synopsys translate_off
defparam \LessThan0~59 .lut_mask = 16'h004D;
defparam \LessThan0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N28
cycloneive_lcell_comb \LessThan0~61 (
// Equation(s):
// \LessThan0~61_cout  = CARRY((Mux1 & (\Selector70~1_combout  & !\LessThan0~59_cout )) # (!Mux1 & ((\Selector70~1_combout ) # (!\LessThan0~59_cout ))))

	.dataa(Mux1),
	.datab(Selector701),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~59_cout ),
	.combout(),
	.cout(\LessThan0~61_cout ));
// synopsys translate_off
defparam \LessThan0~61 .lut_mask = 16'h004D;
defparam \LessThan0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N30
cycloneive_lcell_comb \LessThan0~62 (
// Equation(s):
// \LessThan0~62_combout  = (\Selector69~1_combout  & (\LessThan0~61_cout  & Mux0)) # (!\Selector69~1_combout  & ((\LessThan0~61_cout ) # (Mux0)))

	.dataa(gnd),
	.datab(Selector691),
	.datac(gnd),
	.datad(Mux0),
	.cin(\LessThan0~61_cout ),
	.combout(\LessThan0~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan0~62 .lut_mask = 16'hF330;
defparam \LessThan0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N0
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_cout  = CARRY((!Mux31 & \Selector100~4_combout ))

	.dataa(Mux31),
	.datab(Selector1002),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h0044;
defparam \LessThan1~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N2
cycloneive_lcell_comb \LessThan1~3 (
// Equation(s):
// \LessThan1~3_cout  = CARRY((Mux30 & ((!\LessThan1~1_cout ) # (!\Selector99~2_combout ))) # (!Mux30 & (!\Selector99~2_combout  & !\LessThan1~1_cout )))

	.dataa(Mux30),
	.datab(Selector991),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
// synopsys translate_off
defparam \LessThan1~3 .lut_mask = 16'h002B;
defparam \LessThan1~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N4
cycloneive_lcell_comb \LessThan1~5 (
// Equation(s):
// \LessThan1~5_cout  = CARRY((Mux29 & (\Selector98~2_combout  & !\LessThan1~3_cout )) # (!Mux29 & ((\Selector98~2_combout ) # (!\LessThan1~3_cout ))))

	.dataa(Mux29),
	.datab(Selector981),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
// synopsys translate_off
defparam \LessThan1~5 .lut_mask = 16'h004D;
defparam \LessThan1~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N6
cycloneive_lcell_comb \LessThan1~7 (
// Equation(s):
// \LessThan1~7_cout  = CARRY((Mux28 & ((!\LessThan1~5_cout ) # (!\Selector97~2_combout ))) # (!Mux28 & (!\Selector97~2_combout  & !\LessThan1~5_cout )))

	.dataa(Mux28),
	.datab(Selector971),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
// synopsys translate_off
defparam \LessThan1~7 .lut_mask = 16'h002B;
defparam \LessThan1~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N8
cycloneive_lcell_comb \LessThan1~9 (
// Equation(s):
// \LessThan1~9_cout  = CARRY((Mux27 & (\Selector96~2_combout  & !\LessThan1~7_cout )) # (!Mux27 & ((\Selector96~2_combout ) # (!\LessThan1~7_cout ))))

	.dataa(Mux27),
	.datab(Selector961),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
// synopsys translate_off
defparam \LessThan1~9 .lut_mask = 16'h004D;
defparam \LessThan1~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N10
cycloneive_lcell_comb \LessThan1~11 (
// Equation(s):
// \LessThan1~11_cout  = CARRY((\Selector95~3_combout  & (Mux26 & !\LessThan1~9_cout )) # (!\Selector95~3_combout  & ((Mux26) # (!\LessThan1~9_cout ))))

	.dataa(Selector952),
	.datab(Mux26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
// synopsys translate_off
defparam \LessThan1~11 .lut_mask = 16'h004D;
defparam \LessThan1~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N12
cycloneive_lcell_comb \LessThan1~13 (
// Equation(s):
// \LessThan1~13_cout  = CARRY((Mux25 & (\Selector94~1_combout  & !\LessThan1~11_cout )) # (!Mux25 & ((\Selector94~1_combout ) # (!\LessThan1~11_cout ))))

	.dataa(Mux25),
	.datab(Selector941),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
// synopsys translate_off
defparam \LessThan1~13 .lut_mask = 16'h004D;
defparam \LessThan1~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N14
cycloneive_lcell_comb \LessThan1~15 (
// Equation(s):
// \LessThan1~15_cout  = CARRY((Mux24 & ((!\LessThan1~13_cout ) # (!\Selector93~1_combout ))) # (!Mux24 & (!\Selector93~1_combout  & !\LessThan1~13_cout )))

	.dataa(Mux24),
	.datab(Selector931),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
// synopsys translate_off
defparam \LessThan1~15 .lut_mask = 16'h002B;
defparam \LessThan1~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N16
cycloneive_lcell_comb \LessThan1~17 (
// Equation(s):
// \LessThan1~17_cout  = CARRY((Mux23 & (\Selector92~1_combout  & !\LessThan1~15_cout )) # (!Mux23 & ((\Selector92~1_combout ) # (!\LessThan1~15_cout ))))

	.dataa(Mux23),
	.datab(Selector921),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
// synopsys translate_off
defparam \LessThan1~17 .lut_mask = 16'h004D;
defparam \LessThan1~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N18
cycloneive_lcell_comb \LessThan1~19 (
// Equation(s):
// \LessThan1~19_cout  = CARRY((Mux22 & ((!\LessThan1~17_cout ) # (!\Selector91~1_combout ))) # (!Mux22 & (!\Selector91~1_combout  & !\LessThan1~17_cout )))

	.dataa(Mux22),
	.datab(Selector911),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
// synopsys translate_off
defparam \LessThan1~19 .lut_mask = 16'h002B;
defparam \LessThan1~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N20
cycloneive_lcell_comb \LessThan1~21 (
// Equation(s):
// \LessThan1~21_cout  = CARRY((\Selector90~1_combout  & ((!\LessThan1~19_cout ) # (!Mux21))) # (!\Selector90~1_combout  & (!Mux21 & !\LessThan1~19_cout )))

	.dataa(Selector901),
	.datab(Mux21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
// synopsys translate_off
defparam \LessThan1~21 .lut_mask = 16'h002B;
defparam \LessThan1~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N22
cycloneive_lcell_comb \LessThan1~23 (
// Equation(s):
// \LessThan1~23_cout  = CARRY((Mux20 & ((!\LessThan1~21_cout ) # (!\Selector89~1_combout ))) # (!Mux20 & (!\Selector89~1_combout  & !\LessThan1~21_cout )))

	.dataa(Mux20),
	.datab(Selector891),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
// synopsys translate_off
defparam \LessThan1~23 .lut_mask = 16'h002B;
defparam \LessThan1~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N24
cycloneive_lcell_comb \LessThan1~25 (
// Equation(s):
// \LessThan1~25_cout  = CARRY((Mux19 & (\Selector88~1_combout  & !\LessThan1~23_cout )) # (!Mux19 & ((\Selector88~1_combout ) # (!\LessThan1~23_cout ))))

	.dataa(Mux19),
	.datab(Selector881),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
// synopsys translate_off
defparam \LessThan1~25 .lut_mask = 16'h004D;
defparam \LessThan1~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N26
cycloneive_lcell_comb \LessThan1~27 (
// Equation(s):
// \LessThan1~27_cout  = CARRY((Mux18 & ((!\LessThan1~25_cout ) # (!\Selector87~1_combout ))) # (!Mux18 & (!\Selector87~1_combout  & !\LessThan1~25_cout )))

	.dataa(Mux18),
	.datab(Selector871),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
// synopsys translate_off
defparam \LessThan1~27 .lut_mask = 16'h002B;
defparam \LessThan1~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N28
cycloneive_lcell_comb \LessThan1~29 (
// Equation(s):
// \LessThan1~29_cout  = CARRY((Mux17 & (\Selector86~1_combout  & !\LessThan1~27_cout )) # (!Mux17 & ((\Selector86~1_combout ) # (!\LessThan1~27_cout ))))

	.dataa(Mux17),
	.datab(Selector861),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
// synopsys translate_off
defparam \LessThan1~29 .lut_mask = 16'h004D;
defparam \LessThan1~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N30
cycloneive_lcell_comb \LessThan1~31 (
// Equation(s):
// \LessThan1~31_cout  = CARRY((Mux16 & ((!\LessThan1~29_cout ) # (!\Selector85~1_combout ))) # (!Mux16 & (!\Selector85~1_combout  & !\LessThan1~29_cout )))

	.dataa(Mux16),
	.datab(Selector851),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~29_cout ),
	.combout(),
	.cout(\LessThan1~31_cout ));
// synopsys translate_off
defparam \LessThan1~31 .lut_mask = 16'h002B;
defparam \LessThan1~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N0
cycloneive_lcell_comb \LessThan1~33 (
// Equation(s):
// \LessThan1~33_cout  = CARRY((\Selector84~2_combout  & ((!\LessThan1~31_cout ) # (!Mux15))) # (!\Selector84~2_combout  & (!Mux15 & !\LessThan1~31_cout )))

	.dataa(Selector841),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~31_cout ),
	.combout(),
	.cout(\LessThan1~33_cout ));
// synopsys translate_off
defparam \LessThan1~33 .lut_mask = 16'h002B;
defparam \LessThan1~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N2
cycloneive_lcell_comb \LessThan1~35 (
// Equation(s):
// \LessThan1~35_cout  = CARRY((Mux14 & ((!\LessThan1~33_cout ) # (!\Selector83~1_combout ))) # (!Mux14 & (!\Selector83~1_combout  & !\LessThan1~33_cout )))

	.dataa(Mux14),
	.datab(Selector831),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~33_cout ),
	.combout(),
	.cout(\LessThan1~35_cout ));
// synopsys translate_off
defparam \LessThan1~35 .lut_mask = 16'h002B;
defparam \LessThan1~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N4
cycloneive_lcell_comb \LessThan1~37 (
// Equation(s):
// \LessThan1~37_cout  = CARRY((\Selector82~1_combout  & ((!\LessThan1~35_cout ) # (!Mux13))) # (!\Selector82~1_combout  & (!Mux13 & !\LessThan1~35_cout )))

	.dataa(Selector821),
	.datab(Mux13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~35_cout ),
	.combout(),
	.cout(\LessThan1~37_cout ));
// synopsys translate_off
defparam \LessThan1~37 .lut_mask = 16'h002B;
defparam \LessThan1~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N6
cycloneive_lcell_comb \LessThan1~39 (
// Equation(s):
// \LessThan1~39_cout  = CARRY((Mux12 & ((!\LessThan1~37_cout ) # (!\Selector81~1_combout ))) # (!Mux12 & (!\Selector81~1_combout  & !\LessThan1~37_cout )))

	.dataa(Mux12),
	.datab(Selector811),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~37_cout ),
	.combout(),
	.cout(\LessThan1~39_cout ));
// synopsys translate_off
defparam \LessThan1~39 .lut_mask = 16'h002B;
defparam \LessThan1~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N8
cycloneive_lcell_comb \LessThan1~41 (
// Equation(s):
// \LessThan1~41_cout  = CARRY((Mux11 & (\Selector80~1_combout  & !\LessThan1~39_cout )) # (!Mux11 & ((\Selector80~1_combout ) # (!\LessThan1~39_cout ))))

	.dataa(Mux11),
	.datab(Selector801),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~39_cout ),
	.combout(),
	.cout(\LessThan1~41_cout ));
// synopsys translate_off
defparam \LessThan1~41 .lut_mask = 16'h004D;
defparam \LessThan1~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N10
cycloneive_lcell_comb \LessThan1~43 (
// Equation(s):
// \LessThan1~43_cout  = CARRY((Mux10 & ((!\LessThan1~41_cout ) # (!\Selector79~1_combout ))) # (!Mux10 & (!\Selector79~1_combout  & !\LessThan1~41_cout )))

	.dataa(Mux10),
	.datab(Selector791),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~41_cout ),
	.combout(),
	.cout(\LessThan1~43_cout ));
// synopsys translate_off
defparam \LessThan1~43 .lut_mask = 16'h002B;
defparam \LessThan1~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N12
cycloneive_lcell_comb \LessThan1~45 (
// Equation(s):
// \LessThan1~45_cout  = CARRY((\Selector78~1_combout  & ((!\LessThan1~43_cout ) # (!Mux9))) # (!\Selector78~1_combout  & (!Mux9 & !\LessThan1~43_cout )))

	.dataa(Selector781),
	.datab(Mux9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~43_cout ),
	.combout(),
	.cout(\LessThan1~45_cout ));
// synopsys translate_off
defparam \LessThan1~45 .lut_mask = 16'h002B;
defparam \LessThan1~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N14
cycloneive_lcell_comb \LessThan1~47 (
// Equation(s):
// \LessThan1~47_cout  = CARRY((\Selector77~1_combout  & (Mux8 & !\LessThan1~45_cout )) # (!\Selector77~1_combout  & ((Mux8) # (!\LessThan1~45_cout ))))

	.dataa(Selector771),
	.datab(Mux8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~45_cout ),
	.combout(),
	.cout(\LessThan1~47_cout ));
// synopsys translate_off
defparam \LessThan1~47 .lut_mask = 16'h004D;
defparam \LessThan1~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N16
cycloneive_lcell_comb \LessThan1~49 (
// Equation(s):
// \LessThan1~49_cout  = CARRY((Mux7 & (\Selector76~1_combout  & !\LessThan1~47_cout )) # (!Mux7 & ((\Selector76~1_combout ) # (!\LessThan1~47_cout ))))

	.dataa(Mux7),
	.datab(Selector761),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~47_cout ),
	.combout(),
	.cout(\LessThan1~49_cout ));
// synopsys translate_off
defparam \LessThan1~49 .lut_mask = 16'h004D;
defparam \LessThan1~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N18
cycloneive_lcell_comb \LessThan1~51 (
// Equation(s):
// \LessThan1~51_cout  = CARRY((\Selector75~1_combout  & (Mux6 & !\LessThan1~49_cout )) # (!\Selector75~1_combout  & ((Mux6) # (!\LessThan1~49_cout ))))

	.dataa(Selector751),
	.datab(Mux6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~49_cout ),
	.combout(),
	.cout(\LessThan1~51_cout ));
// synopsys translate_off
defparam \LessThan1~51 .lut_mask = 16'h004D;
defparam \LessThan1~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N20
cycloneive_lcell_comb \LessThan1~53 (
// Equation(s):
// \LessThan1~53_cout  = CARRY((Mux5 & (\Selector74~1_combout  & !\LessThan1~51_cout )) # (!Mux5 & ((\Selector74~1_combout ) # (!\LessThan1~51_cout ))))

	.dataa(Mux5),
	.datab(Selector741),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~51_cout ),
	.combout(),
	.cout(\LessThan1~53_cout ));
// synopsys translate_off
defparam \LessThan1~53 .lut_mask = 16'h004D;
defparam \LessThan1~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N22
cycloneive_lcell_comb \LessThan1~55 (
// Equation(s):
// \LessThan1~55_cout  = CARRY((\Selector73~1_combout  & (Mux4 & !\LessThan1~53_cout )) # (!\Selector73~1_combout  & ((Mux4) # (!\LessThan1~53_cout ))))

	.dataa(Selector731),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~53_cout ),
	.combout(),
	.cout(\LessThan1~55_cout ));
// synopsys translate_off
defparam \LessThan1~55 .lut_mask = 16'h004D;
defparam \LessThan1~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N24
cycloneive_lcell_comb \LessThan1~57 (
// Equation(s):
// \LessThan1~57_cout  = CARRY((\Selector72~1_combout  & ((!\LessThan1~55_cout ) # (!Mux3))) # (!\Selector72~1_combout  & (!Mux3 & !\LessThan1~55_cout )))

	.dataa(Selector721),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~55_cout ),
	.combout(),
	.cout(\LessThan1~57_cout ));
// synopsys translate_off
defparam \LessThan1~57 .lut_mask = 16'h002B;
defparam \LessThan1~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N26
cycloneive_lcell_comb \LessThan1~59 (
// Equation(s):
// \LessThan1~59_cout  = CARRY((\Selector71~1_combout  & (Mux2 & !\LessThan1~57_cout )) # (!\Selector71~1_combout  & ((Mux2) # (!\LessThan1~57_cout ))))

	.dataa(Selector711),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~57_cout ),
	.combout(),
	.cout(\LessThan1~59_cout ));
// synopsys translate_off
defparam \LessThan1~59 .lut_mask = 16'h004D;
defparam \LessThan1~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N28
cycloneive_lcell_comb \LessThan1~61 (
// Equation(s):
// \LessThan1~61_cout  = CARRY((Mux1 & (\Selector70~1_combout  & !\LessThan1~59_cout )) # (!Mux1 & ((\Selector70~1_combout ) # (!\LessThan1~59_cout ))))

	.dataa(Mux1),
	.datab(Selector701),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~59_cout ),
	.combout(),
	.cout(\LessThan1~61_cout ));
// synopsys translate_off
defparam \LessThan1~61 .lut_mask = 16'h004D;
defparam \LessThan1~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N30
cycloneive_lcell_comb \LessThan1~62 (
// Equation(s):
// \LessThan1~62_combout  = (\Selector69~1_combout  & ((\LessThan1~61_cout ) # (!Mux0))) # (!\Selector69~1_combout  & (\LessThan1~61_cout  & !Mux0))

	.dataa(gnd),
	.datab(Selector691),
	.datac(gnd),
	.datad(Mux0),
	.cin(\LessThan1~61_cout ),
	.combout(\LessThan1~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~62 .lut_mask = 16'hC0FC;
defparam \LessThan1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N0
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (\Mux31~1_combout  & ((Selector3 & ((\LessThan1~62_combout ))) # (!Selector3 & (\LessThan0~62_combout ))))

	.dataa(\Mux31~1_combout ),
	.datab(Selector3),
	.datac(\LessThan0~62_combout ),
	.datad(\LessThan1~62_combout ),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hA820;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N2
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (Mux31 & (Selector2 $ (((Selector3) # (\Selector100~4_combout ))))) # (!Mux31 & ((Selector2 & (Selector3 $ (\Selector100~4_combout ))) # (!Selector2 & (Selector3 & \Selector100~4_combout ))))

	.dataa(Mux31),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector1002),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'h3668;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N4
cycloneive_lcell_comb \Equal0~6 (
// Equation(s):
// \Equal0~6_combout  = (!Mux103 & (!Mux93 & ((!\Mux31~3_combout ) # (!Mux311))))

	.dataa(Mux311),
	.datab(Mux103),
	.datac(\Mux31~3_combout ),
	.datad(Mux93),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~6 .lut_mask = 16'h0013;
defparam \Equal0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N4
cycloneive_lcell_comb \Equal0~3 (
// Equation(s):
// \Equal0~3_combout  = (!Mux223 & (!Mux233 & (!Mux213 & !Mux203)))

	.dataa(Mux223),
	.datab(Mux233),
	.datac(Mux213),
	.datad(Mux203),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~3 .lut_mask = 16'h0001;
defparam \Equal0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N2
cycloneive_lcell_comb \Equal0~4 (
// Equation(s):
// \Equal0~4_combout  = (!Mux173 & (!Mux193 & (!Mux163 & !Mux183)))

	.dataa(Mux173),
	.datab(Mux193),
	.datac(Mux163),
	.datad(Mux183),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~4 .lut_mask = 16'h0001;
defparam \Equal0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N24
cycloneive_lcell_comb \Equal0~5 (
// Equation(s):
// \Equal0~5_combout  = (!Mux291 & (!Mux281 & (\Equal0~3_combout  & \Equal0~4_combout )))

	.dataa(Mux291),
	.datab(Mux281),
	.datac(\Equal0~3_combout ),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~5 .lut_mask = 16'h1000;
defparam \Equal0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N20
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (\Selector100~4_combout  & (Selector3 & ((Mux30)))) # (!\Selector100~4_combout  & (((Mux31))))

	.dataa(Selector1002),
	.datab(Selector3),
	.datac(Mux31),
	.datad(Mux30),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hD850;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N14
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (\Selector99~2_combout  & (Selector3 & (\ShiftRight0~90_combout ))) # (!\Selector99~2_combout  & (((\Mux31~4_combout ))))

	.dataa(Selector991),
	.datab(Selector3),
	.datac(\ShiftRight0~90_combout ),
	.datad(\Mux31~4_combout ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hD580;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N24
cycloneive_lcell_comb \ShiftRight0~67 (
// Equation(s):
// \ShiftRight0~67_combout  = (\Selector99~2_combout  & ((\Selector100~4_combout  & (Mux24)) # (!\Selector100~4_combout  & ((Mux25)))))

	.dataa(Mux24),
	.datab(Selector991),
	.datac(Mux25),
	.datad(Selector1002),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~67 .lut_mask = 16'h88C0;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N0
cycloneive_lcell_comb \ShiftRight0~69 (
// Equation(s):
// \ShiftRight0~69_combout  = (\ShiftRight0~67_combout ) # ((!\Selector99~2_combout  & \ShiftRight0~68_combout ))

	.dataa(gnd),
	.datab(Selector991),
	.datac(\ShiftRight0~68_combout ),
	.datad(\ShiftRight0~67_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~69 .lut_mask = 16'hFF30;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N22
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (\Selector98~2_combout  & (Selector3 & ((\ShiftRight0~69_combout )))) # (!\Selector98~2_combout  & (((\Mux31~5_combout ))))

	.dataa(Selector3),
	.datab(Selector981),
	.datac(\Mux31~5_combout ),
	.datad(\ShiftRight0~69_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hB830;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N16
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (\Selector97~2_combout  & (Selector3 & ((\ShiftRight0~83_combout )))) # (!\Selector97~2_combout  & (((\Mux31~6_combout ))))

	.dataa(Selector3),
	.datab(Selector971),
	.datac(\Mux31~6_combout ),
	.datad(\ShiftRight0~83_combout ),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hB830;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N14
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (\Mux0~4_combout  & (!Selector2 & \Mux31~7_combout ))

	.dataa(\Mux0~4_combout ),
	.datab(gnd),
	.datac(Selector2),
	.datad(\Mux31~7_combout ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'h0A00;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N8
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// \Mux31~9_combout  = (\Selector96~2_combout  & (\Mux6~17_combout  & (!\ShiftLeft0~32_combout  & \ShiftRight0~102_combout )))

	.dataa(Selector961),
	.datab(\Mux6~17_combout ),
	.datac(\ShiftLeft0~32_combout ),
	.datad(\ShiftRight0~102_combout ),
	.cin(gnd),
	.combout(\Mux31~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'h0800;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N6
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (\Mux31~9_combout ) # ((Selector2 & \Add0~33_combout ))

	.dataa(gnd),
	.datab(Selector2),
	.datac(\Mux31~9_combout ),
	.datad(\Add0~33_combout ),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hFCF0;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N0
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (!Selector0 & (!Selector1 & ((\Mux31~8_combout ) # (\Mux31~10_combout ))))

	.dataa(Selector0),
	.datab(Selector1),
	.datac(\Mux31~8_combout ),
	.datad(\Mux31~10_combout ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'h1110;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N30
cycloneive_lcell_comb \Equal0~7 (
// Equation(s):
// \Equal0~7_combout  = (!Mux123 & (!Mux153 & (!Mux143 & !Mux133)))

	.dataa(Mux123),
	.datab(Mux153),
	.datac(Mux143),
	.datad(Mux133),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~7 .lut_mask = 16'h0001;
defparam \Equal0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N2
cycloneive_lcell_comb \Equal0~8 (
// Equation(s):
// \Equal0~8_combout  = (!Mux301 & (!\Mux31~11_combout  & (!Mux115 & \Equal0~7_combout )))

	.dataa(Mux301),
	.datab(\Mux31~11_combout ),
	.datac(Mux115),
	.datad(\Equal0~7_combout ),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~8 .lut_mask = 16'h0100;
defparam \Equal0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N20
cycloneive_lcell_comb \Equal0~9 (
// Equation(s):
// \Equal0~9_combout  = (\Equal0~6_combout  & (!Mux81 & (\Equal0~5_combout  & \Equal0~8_combout )))

	.dataa(\Equal0~6_combout ),
	.datab(Mux81),
	.datac(\Equal0~5_combout ),
	.datad(\Equal0~8_combout ),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~9 .lut_mask = 16'h2000;
defparam \Equal0~9 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module control_unit (
	always1,
	ccifiwait_0,
	dcifimemload_26,
	dcifimemload_27,
	dcifimemload_28,
	dcifimemload_29,
	dcifimemload_30,
	dcifimemload_31,
	dcifihit,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_0,
	dcifimemload_1,
	Selector5,
	nxtwen,
	WideOr3,
	cuifALUSrc_1,
	Decoder1,
	WideOr13,
	Selector3,
	Selector0,
	Selector1,
	Selector2,
	Equal0,
	Equal01,
	Selector6,
	cuifRegSel_0,
	cuifRegSel_1,
	Decoder11,
	Selector4,
	Selector41,
	Selector42,
	Mux1,
	cuifRegSel_11,
	devpor,
	devclrn,
	devoe);
input 	always1;
input 	ccifiwait_0;
input 	dcifimemload_26;
input 	dcifimemload_27;
input 	dcifimemload_28;
input 	dcifimemload_29;
input 	dcifimemload_30;
input 	dcifimemload_31;
input 	dcifihit;
input 	dcifimemload_3;
input 	dcifimemload_4;
input 	dcifimemload_2;
input 	dcifimemload_5;
input 	dcifimemload_0;
input 	dcifimemload_1;
output 	Selector5;
input 	nxtwen;
output 	WideOr3;
output 	cuifALUSrc_1;
output 	Decoder1;
output 	WideOr13;
output 	Selector3;
output 	Selector0;
output 	Selector1;
output 	Selector2;
input 	Equal0;
input 	Equal01;
output 	Selector6;
output 	cuifRegSel_0;
output 	cuifRegSel_1;
output 	Decoder11;
output 	Selector4;
output 	Selector41;
output 	Selector42;
input 	Mux1;
output 	cuifRegSel_11;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Decoder1~0_combout ;
wire \Decoder0~0_combout ;
wire \cuif.ALUSrc[1]~4_combout ;
wire \cuif.ALUSrc[1]~6_combout ;
wire \Selector5~3_combout ;
wire \WideOr3~0_combout ;
wire \Selector3~0_combout ;
wire \Selector3~1_combout ;
wire \Selector1~0_combout ;
wire \Selector3~2_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \Selector1~2_combout ;
wire \Selector1~1_combout ;
wire \WideOr1~0_combout ;
wire \Selector2~0_combout ;
wire \Selector6~0_combout ;
wire \cuif.RegSel[0]~2_combout ;
wire \Decoder0~1_combout ;
wire \Selector4~1_combout ;


// Location: LCCOMB_X55_Y40_N26
cycloneive_lcell_comb \Selector5~2 (
// Equation(s):
// Selector5 = (\Selector5~3_combout ) # ((\Decoder1~0_combout  & (!dcifimemload_28 & dcifimemload_27)))

	.dataa(\Decoder1~0_combout ),
	.datab(\Selector5~3_combout ),
	.datac(dcifimemload_28),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(Selector5),
	.cout());
// synopsys translate_off
defparam \Selector5~2 .lut_mask = 16'hCECC;
defparam \Selector5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N24
cycloneive_lcell_comb \WideOr3~1 (
// Equation(s):
// WideOr3 = (!dcifimemload_30 & ((dcifimemload_29 & (!\WideOr3~0_combout )) # (!dcifimemload_29 & ((nxtwen)))))

	.dataa(\WideOr3~0_combout ),
	.datab(dcifimemload_30),
	.datac(dcifimemload_29),
	.datad(nxtwen),
	.cin(gnd),
	.combout(WideOr3),
	.cout());
// synopsys translate_off
defparam \WideOr3~1 .lut_mask = 16'h1310;
defparam \WideOr3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N28
cycloneive_lcell_comb \cuif.ALUSrc[1]~5 (
// Equation(s):
// cuifALUSrc_1 = (!dcifimemload_3 & (\Decoder0~0_combout  & (\Decoder1~0_combout  & \cuif.ALUSrc[1]~4_combout )))

	.dataa(dcifimemload_3),
	.datab(\Decoder0~0_combout ),
	.datac(\Decoder1~0_combout ),
	.datad(\cuif.ALUSrc[1]~4_combout ),
	.cin(gnd),
	.combout(cuifALUSrc_1),
	.cout());
// synopsys translate_off
defparam \cuif.ALUSrc[1]~5 .lut_mask = 16'h4000;
defparam \cuif.ALUSrc[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N4
cycloneive_lcell_comb \Decoder1~1 (
// Equation(s):
// Decoder1 = (!dcifimemload_30 & !dcifimemload_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(dcifimemload_30),
	.datad(dcifimemload_31),
	.cin(gnd),
	.combout(Decoder1),
	.cout());
// synopsys translate_off
defparam \Decoder1~1 .lut_mask = 16'h000F;
defparam \Decoder1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N6
cycloneive_lcell_comb \WideOr13~0 (
// Equation(s):
// WideOr13 = (!dcifimemload_28 & (dcifimemload_29 & ((!dcifimemload_27) # (!dcifimemload_26))))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_26),
	.datac(dcifimemload_29),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(WideOr13),
	.cout());
// synopsys translate_off
defparam \WideOr13~0 .lut_mask = 16'h1050;
defparam \WideOr13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N2
cycloneive_lcell_comb \Selector3~3 (
// Equation(s):
// Selector3 = (\Selector3~2_combout ) # ((Decoder1 & (\Selector3~0_combout  & !\cuif.ALUSrc[1]~6_combout )))

	.dataa(Decoder1),
	.datab(\Selector3~0_combout ),
	.datac(\cuif.ALUSrc[1]~6_combout ),
	.datad(\Selector3~2_combout ),
	.cin(gnd),
	.combout(Selector3),
	.cout());
// synopsys translate_off
defparam \Selector3~3 .lut_mask = 16'hFF08;
defparam \Selector3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N16
cycloneive_lcell_comb \Selector0~2 (
// Equation(s):
// Selector0 = (\Selector0~0_combout ) # ((!dcifimemload_4 & (\Selector0~1_combout  & \cuif.ALUSrc[1]~6_combout )))

	.dataa(dcifimemload_4),
	.datab(\Selector0~0_combout ),
	.datac(\Selector0~1_combout ),
	.datad(\cuif.ALUSrc[1]~6_combout ),
	.cin(gnd),
	.combout(Selector0),
	.cout());
// synopsys translate_off
defparam \Selector0~2 .lut_mask = 16'hDCCC;
defparam \Selector0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N6
cycloneive_lcell_comb \Selector1~3 (
// Equation(s):
// Selector1 = (\Selector1~1_combout ) # ((\Selector1~2_combout  & ((!dcifimemload_27) # (!dcifimemload_26))))

	.dataa(dcifimemload_26),
	.datab(\Selector1~2_combout ),
	.datac(dcifimemload_27),
	.datad(\Selector1~1_combout ),
	.cin(gnd),
	.combout(Selector1),
	.cout());
// synopsys translate_off
defparam \Selector1~3 .lut_mask = 16'hFF4C;
defparam \Selector1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N12
cycloneive_lcell_comb \Selector2~1 (
// Equation(s):
// Selector2 = (\Selector2~0_combout  & ((dcifimemload_3) # ((\WideOr1~0_combout ) # (!\Selector1~0_combout ))))

	.dataa(dcifimemload_3),
	.datab(\Selector1~0_combout ),
	.datac(\WideOr1~0_combout ),
	.datad(\Selector2~0_combout ),
	.cin(gnd),
	.combout(Selector2),
	.cout());
// synopsys translate_off
defparam \Selector2~1 .lut_mask = 16'hFB00;
defparam \Selector2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N30
cycloneive_lcell_comb \Selector6~1 (
// Equation(s):
// Selector6 = (\Decoder1~0_combout  & ((dcifimemload_28 & (!dcifimemload_27 & \Selector6~0_combout )) # (!dcifimemload_28 & (dcifimemload_27))))

	.dataa(\Decoder1~0_combout ),
	.datab(dcifimemload_28),
	.datac(dcifimemload_27),
	.datad(\Selector6~0_combout ),
	.cin(gnd),
	.combout(Selector6),
	.cout());
// synopsys translate_off
defparam \Selector6~1 .lut_mask = 16'h2820;
defparam \Selector6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N14
cycloneive_lcell_comb \cuif.RegSel[0]~3 (
// Equation(s):
// cuifRegSel_0 = (!dcifimemload_30 & (dcifimemload_27 & \cuif.RegSel[0]~2_combout ))

	.dataa(dcifimemload_30),
	.datab(dcifimemload_27),
	.datac(gnd),
	.datad(\cuif.RegSel[0]~2_combout ),
	.cin(gnd),
	.combout(cuifRegSel_0),
	.cout());
// synopsys translate_off
defparam \cuif.RegSel[0]~3 .lut_mask = 16'h4400;
defparam \cuif.RegSel[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N18
cycloneive_lcell_comb \cuif.RegSel[1]~4 (
// Equation(s):
// cuifRegSel_1 = (dcifimemload_27 & (dcifimemload_26 & (dcifimemload_28 $ (!dcifimemload_29))))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_29),
	.datac(dcifimemload_27),
	.datad(dcifimemload_26),
	.cin(gnd),
	.combout(cuifRegSel_1),
	.cout());
// synopsys translate_off
defparam \cuif.RegSel[1]~4 .lut_mask = 16'h9000;
defparam \cuif.RegSel[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N8
cycloneive_lcell_comb \Decoder1~2 (
// Equation(s):
// Decoder11 = (!dcifimemload_28 & (dcifimemload_26 & dcifimemload_27))

	.dataa(dcifimemload_28),
	.datab(gnd),
	.datac(dcifimemload_26),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(Decoder11),
	.cout());
// synopsys translate_off
defparam \Decoder1~2 .lut_mask = 16'h5000;
defparam \Decoder1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N12
cycloneive_lcell_comb \Selector4~0 (
// Equation(s):
// Selector4 = (always1 & (!ccifiwait_0 & (!dcifimemload_29 & nxtwen)))

	.dataa(always1),
	.datab(ccifiwait_0),
	.datac(dcifimemload_29),
	.datad(nxtwen),
	.cin(gnd),
	.combout(Selector4),
	.cout());
// synopsys translate_off
defparam \Selector4~0 .lut_mask = 16'h0200;
defparam \Selector4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N28
cycloneive_lcell_comb \Selector4~2 (
// Equation(s):
// Selector41 = (dcifihit & (!dcifimemload_31 & ((dcifimemload_29) # (\Selector4~1_combout ))))

	.dataa(dcifihit),
	.datab(dcifimemload_29),
	.datac(\Selector4~1_combout ),
	.datad(dcifimemload_31),
	.cin(gnd),
	.combout(Selector41),
	.cout());
// synopsys translate_off
defparam \Selector4~2 .lut_mask = 16'h00A8;
defparam \Selector4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N4
cycloneive_lcell_comb \Selector4~3 (
// Equation(s):
// Selector42 = (!dcifimemload_30 & ((Selector4) # (Selector41)))

	.dataa(Selector4),
	.datab(gnd),
	.datac(dcifimemload_30),
	.datad(Selector41),
	.cin(gnd),
	.combout(Selector42),
	.cout());
// synopsys translate_off
defparam \Selector4~3 .lut_mask = 16'h0F0A;
defparam \Selector4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N24
cycloneive_lcell_comb \cuif.RegSel[1]~5 (
// Equation(s):
// cuifRegSel_11 = (!dcifimemload_31 & (cuifRegSel_1 & !dcifimemload_30))

	.dataa(dcifimemload_31),
	.datab(gnd),
	.datac(cuifRegSel_1),
	.datad(dcifimemload_30),
	.cin(gnd),
	.combout(cuifRegSel_11),
	.cout());
// synopsys translate_off
defparam \cuif.RegSel[1]~5 .lut_mask = 16'h0050;
defparam \cuif.RegSel[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N22
cycloneive_lcell_comb \Decoder1~0 (
// Equation(s):
// \Decoder1~0_combout  = (!dcifimemload_31 & (!dcifimemload_29 & !dcifimemload_30))

	.dataa(gnd),
	.datab(dcifimemload_31),
	.datac(dcifimemload_29),
	.datad(dcifimemload_30),
	.cin(gnd),
	.combout(\Decoder1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder1~0 .lut_mask = 16'h0003;
defparam \Decoder1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N16
cycloneive_lcell_comb \Decoder0~0 (
// Equation(s):
// \Decoder0~0_combout  = (!dcifimemload_2 & (!dcifimemload_5 & (!dcifimemload_4 & !dcifimemload_0)))

	.dataa(dcifimemload_2),
	.datab(dcifimemload_5),
	.datac(dcifimemload_4),
	.datad(dcifimemload_0),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~0 .lut_mask = 16'h0001;
defparam \Decoder0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N0
cycloneive_lcell_comb \cuif.ALUSrc[1]~4 (
// Equation(s):
// \cuif.ALUSrc[1]~4_combout  = (!dcifimemload_28 & (!dcifimemload_27 & !dcifimemload_26))

	.dataa(gnd),
	.datab(dcifimemload_28),
	.datac(dcifimemload_27),
	.datad(dcifimemload_26),
	.cin(gnd),
	.combout(\cuif.ALUSrc[1]~4_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUSrc[1]~4 .lut_mask = 16'h0003;
defparam \cuif.ALUSrc[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N10
cycloneive_lcell_comb \cuif.ALUSrc[1]~6 (
// Equation(s):
// \cuif.ALUSrc[1]~6_combout  = (!dcifimemload_31 & (!dcifimemload_30 & (!dcifimemload_29 & \cuif.ALUSrc[1]~4_combout )))

	.dataa(dcifimemload_31),
	.datab(dcifimemload_30),
	.datac(dcifimemload_29),
	.datad(\cuif.ALUSrc[1]~4_combout ),
	.cin(gnd),
	.combout(\cuif.ALUSrc[1]~6_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUSrc[1]~6 .lut_mask = 16'h0100;
defparam \cuif.ALUSrc[1]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N14
cycloneive_lcell_comb \Selector5~3 (
// Equation(s):
// \Selector5~3_combout  = (dcifimemload_3 & (\Decoder0~0_combout  & (!dcifimemload_1 & \cuif.ALUSrc[1]~6_combout )))

	.dataa(dcifimemload_3),
	.datab(\Decoder0~0_combout ),
	.datac(dcifimemload_1),
	.datad(\cuif.ALUSrc[1]~6_combout ),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~3 .lut_mask = 16'h0800;
defparam \Selector5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N26
cycloneive_lcell_comb \WideOr3~0 (
// Equation(s):
// \WideOr3~0_combout  = (dcifimemload_26 & ((dcifimemload_27 & ((dcifimemload_28))) # (!dcifimemload_27 & (dcifimemload_31)))) # (!dcifimemload_26 & (((dcifimemload_31))))

	.dataa(dcifimemload_26),
	.datab(dcifimemload_27),
	.datac(dcifimemload_31),
	.datad(dcifimemload_28),
	.cin(gnd),
	.combout(\WideOr3~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr3~0 .lut_mask = 16'hF870;
defparam \WideOr3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N16
cycloneive_lcell_comb \Selector3~0 (
// Equation(s):
// \Selector3~0_combout  = (dcifimemload_29 & (dcifimemload_26 & (dcifimemload_28 $ (dcifimemload_27)))) # (!dcifimemload_29 & (dcifimemload_28 & ((!dcifimemload_27))))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_26),
	.datac(dcifimemload_27),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~0 .lut_mask = 16'h480A;
defparam \Selector3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N26
cycloneive_lcell_comb \Selector3~1 (
// Equation(s):
// \Selector3~1_combout  = (dcifimemload_3 & (!dcifimemload_2 & ((!dcifimemload_0) # (!dcifimemload_5)))) # (!dcifimemload_3 & (dcifimemload_0 & (dcifimemload_5 $ (!dcifimemload_2))))

	.dataa(dcifimemload_3),
	.datab(dcifimemload_5),
	.datac(dcifimemload_2),
	.datad(dcifimemload_0),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~1 .lut_mask = 16'h430A;
defparam \Selector3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N28
cycloneive_lcell_comb \Selector1~0 (
// Equation(s):
// \Selector1~0_combout  = (\cuif.ALUSrc[1]~4_combout  & (\Decoder1~0_combout  & !dcifimemload_4))

	.dataa(gnd),
	.datab(\cuif.ALUSrc[1]~4_combout ),
	.datac(\Decoder1~0_combout ),
	.datad(dcifimemload_4),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~0 .lut_mask = 16'h00C0;
defparam \Selector1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N12
cycloneive_lcell_comb \Selector3~2 (
// Equation(s):
// \Selector3~2_combout  = (\Selector1~0_combout  & ((dcifimemload_2 & ((\Selector3~1_combout ))) # (!dcifimemload_2 & (dcifimemload_1 & !\Selector3~1_combout ))))

	.dataa(dcifimemload_2),
	.datab(dcifimemload_1),
	.datac(\Selector3~1_combout ),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~2 .lut_mask = 16'hA400;
defparam \Selector3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N24
cycloneive_lcell_comb \Selector0~0 (
// Equation(s):
// \Selector0~0_combout  = (!dcifimemload_28 & (dcifimemload_27 & (Decoder1 & dcifimemload_29)))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_27),
	.datac(Decoder1),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~0 .lut_mask = 16'h4000;
defparam \Selector0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N26
cycloneive_lcell_comb \Selector0~1 (
// Equation(s):
// \Selector0~1_combout  = (dcifimemload_3 & (dcifimemload_5 & (dcifimemload_1 & !dcifimemload_2)))

	.dataa(dcifimemload_3),
	.datab(dcifimemload_5),
	.datac(dcifimemload_1),
	.datad(dcifimemload_2),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~1 .lut_mask = 16'h0080;
defparam \Selector0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N0
cycloneive_lcell_comb \Selector1~2 (
// Equation(s):
// \Selector1~2_combout  = (dcifimemload_28 & (dcifimemload_29 & (!dcifimemload_30 & !dcifimemload_31)))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_29),
	.datac(dcifimemload_30),
	.datad(dcifimemload_31),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~2 .lut_mask = 16'h0008;
defparam \Selector1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N2
cycloneive_lcell_comb \Selector1~1 (
// Equation(s):
// \Selector1~1_combout  = (dcifimemload_5 & (!dcifimemload_3 & (\Selector1~0_combout  & dcifimemload_2)))

	.dataa(dcifimemload_5),
	.datab(dcifimemload_3),
	.datac(\Selector1~0_combout ),
	.datad(dcifimemload_2),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~1 .lut_mask = 16'h2000;
defparam \Selector1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N22
cycloneive_lcell_comb \WideOr1~0 (
// Equation(s):
// \WideOr1~0_combout  = (dcifimemload_2 & (((dcifimemload_1) # (!dcifimemload_5)))) # (!dcifimemload_2 & ((dcifimemload_0) # ((dcifimemload_5))))

	.dataa(dcifimemload_0),
	.datab(dcifimemload_2),
	.datac(dcifimemload_1),
	.datad(dcifimemload_5),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~0 .lut_mask = 16'hF3EE;
defparam \WideOr1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N22
cycloneive_lcell_comb \Selector2~0 (
// Equation(s):
// \Selector2~0_combout  = ((dcifimemload_27) # ((!dcifimemload_29) # (!Decoder1))) # (!dcifimemload_28)

	.dataa(dcifimemload_28),
	.datab(dcifimemload_27),
	.datac(Decoder1),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~0 .lut_mask = 16'hDFFF;
defparam \Selector2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N24
cycloneive_lcell_comb \Selector6~0 (
// Equation(s):
// \Selector6~0_combout  = dcifimemload_26 $ (((!Mux114 & (Equal0 & Equal01))))

	.dataa(dcifimemload_26),
	.datab(Mux1),
	.datac(Equal0),
	.datad(Equal01),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~0 .lut_mask = 16'h9AAA;
defparam \Selector6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N24
cycloneive_lcell_comb \cuif.RegSel[0]~2 (
// Equation(s):
// \cuif.RegSel[0]~2_combout  = (dcifimemload_26 & ((dcifimemload_28 & (dcifimemload_29 & !dcifimemload_31)) # (!dcifimemload_28 & (!dcifimemload_29 & dcifimemload_31))))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_26),
	.datac(dcifimemload_29),
	.datad(dcifimemload_31),
	.cin(gnd),
	.combout(\cuif.RegSel[0]~2_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.RegSel[0]~2 .lut_mask = 16'h0480;
defparam \cuif.RegSel[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N28
cycloneive_lcell_comb \Decoder0~1 (
// Equation(s):
// \Decoder0~1_combout  = (dcifimemload_3 & (\Decoder0~0_combout  & !dcifimemload_1))

	.dataa(dcifimemload_3),
	.datab(gnd),
	.datac(\Decoder0~0_combout ),
	.datad(dcifimemload_1),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~1 .lut_mask = 16'h00A0;
defparam \Decoder0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N26
cycloneive_lcell_comb \Selector4~1 (
// Equation(s):
// \Selector4~1_combout  = (!dcifimemload_28 & ((dcifimemload_26 & (dcifimemload_27)) # (!dcifimemload_26 & (!dcifimemload_27 & !\Decoder0~1_combout ))))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_26),
	.datac(dcifimemload_27),
	.datad(\Decoder0~1_combout ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~1 .lut_mask = 16'h4041;
defparam \Selector4~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module register_file (
	Add1,
	Add11,
	Add12,
	Add13,
	Add14,
	Add15,
	Add16,
	Add17,
	Add18,
	Add19,
	Add110,
	Add111,
	Add112,
	Add113,
	Add114,
	Add115,
	Add116,
	Add117,
	PC_1,
	PC_0,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	dcifimemload_30,
	dcifimemload_31,
	dcifimemload_19,
	dcifimemload_18,
	dcifimemload_16,
	dcifimemload_17,
	Mux63,
	Mux631,
	dcifimemload_24,
	dcifimemload_23,
	dcifimemload_21,
	dcifimemload_22,
	dcifimemload_25,
	Mux30,
	Mux33,
	Mux331,
	Mux1,
	Mux34,
	Mux341,
	Mux2,
	Mux35,
	Mux351,
	Mux3,
	Mux36,
	Mux361,
	Mux4,
	Mux37,
	Mux371,
	Mux5,
	Mux38,
	Mux381,
	Mux6,
	Mux39,
	Mux391,
	Mux7,
	Mux40,
	Mux401,
	Mux8,
	Mux41,
	Mux411,
	Mux9,
	Mux42,
	Mux421,
	Mux10,
	Mux43,
	Mux431,
	Mux11,
	Mux44,
	Mux441,
	Mux12,
	Mux45,
	Mux451,
	Mux13,
	Mux46,
	Mux461,
	Mux14,
	Mux47,
	Mux471,
	Mux15,
	Mux48,
	Mux481,
	Mux16,
	Mux49,
	Mux491,
	Mux17,
	Mux50,
	Mux501,
	Mux18,
	Mux51,
	Mux511,
	Mux19,
	Mux52,
	Mux521,
	dcifimemload_11,
	Mux20,
	Mux53,
	Mux531,
	dcifimemload_10,
	Mux21,
	Mux54,
	Mux541,
	dcifimemload_9,
	Mux22,
	Mux55,
	Mux551,
	dcifimemload_8,
	Mux23,
	Mux56,
	Mux561,
	Mux24,
	Mux57,
	Mux571,
	Mux25,
	Mux58,
	Mux581,
	Mux26,
	Mux59,
	Mux591,
	Mux27,
	Mux60,
	Mux601,
	Mux28,
	Mux61,
	Mux611,
	Mux29,
	Mux62,
	Mux621,
	Mux31,
	Mux32,
	Mux321,
	Mux0,
	Selector0,
	Mux241,
	Mux251,
	Mux261,
	Mux271,
	Mux410,
	Mux510,
	Mux64,
	Mux71,
	Mux291,
	Mux281,
	Mux301,
	Mux311,
	cuifRegSel_0,
	cuifRegSel_1,
	Selector68,
	Selector67,
	Selector64,
	Selector66,
	Selector65,
	Selector4,
	Selector41,
	Selector42,
	Selector1,
	Selector2,
	Selector3,
	Selector8,
	Selector9,
	Selector10,
	Selector11,
	Selector12,
	Selector13,
	Selector14,
	Selector15,
	Selector01,
	Mux231,
	Mux221,
	Mux211,
	Mux201,
	Mux191,
	Mux181,
	Mux171,
	Mux161,
	cuifRegSel_11,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	Add1;
input 	Add11;
input 	Add12;
input 	Add13;
input 	Add14;
input 	Add15;
input 	Add16;
input 	Add17;
input 	Add18;
input 	Add19;
input 	Add110;
input 	Add111;
input 	Add112;
input 	Add113;
input 	Add114;
input 	Add115;
input 	Add116;
input 	Add117;
input 	PC_1;
input 	PC_0;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	dcifimemload_30;
input 	dcifimemload_31;
input 	dcifimemload_19;
input 	dcifimemload_18;
input 	dcifimemload_16;
input 	dcifimemload_17;
output 	Mux63;
output 	Mux631;
input 	dcifimemload_24;
input 	dcifimemload_23;
input 	dcifimemload_21;
input 	dcifimemload_22;
input 	dcifimemload_25;
output 	Mux30;
output 	Mux33;
output 	Mux331;
output 	Mux1;
output 	Mux34;
output 	Mux341;
output 	Mux2;
output 	Mux35;
output 	Mux351;
output 	Mux3;
output 	Mux36;
output 	Mux361;
output 	Mux4;
output 	Mux37;
output 	Mux371;
output 	Mux5;
output 	Mux38;
output 	Mux381;
output 	Mux6;
output 	Mux39;
output 	Mux391;
output 	Mux7;
output 	Mux40;
output 	Mux401;
output 	Mux8;
output 	Mux41;
output 	Mux411;
output 	Mux9;
output 	Mux42;
output 	Mux421;
output 	Mux10;
output 	Mux43;
output 	Mux431;
output 	Mux11;
output 	Mux44;
output 	Mux441;
output 	Mux12;
output 	Mux45;
output 	Mux451;
output 	Mux13;
output 	Mux46;
output 	Mux461;
output 	Mux14;
output 	Mux47;
output 	Mux471;
output 	Mux15;
output 	Mux48;
output 	Mux481;
output 	Mux16;
output 	Mux49;
output 	Mux491;
output 	Mux17;
output 	Mux50;
output 	Mux501;
output 	Mux18;
output 	Mux51;
output 	Mux511;
output 	Mux19;
output 	Mux52;
output 	Mux521;
input 	dcifimemload_11;
output 	Mux20;
output 	Mux53;
output 	Mux531;
input 	dcifimemload_10;
output 	Mux21;
output 	Mux54;
output 	Mux541;
input 	dcifimemload_9;
output 	Mux22;
output 	Mux55;
output 	Mux551;
input 	dcifimemload_8;
output 	Mux23;
output 	Mux56;
output 	Mux561;
output 	Mux24;
output 	Mux57;
output 	Mux571;
output 	Mux25;
output 	Mux58;
output 	Mux581;
output 	Mux26;
output 	Mux59;
output 	Mux591;
output 	Mux27;
output 	Mux60;
output 	Mux601;
output 	Mux28;
output 	Mux61;
output 	Mux611;
output 	Mux29;
output 	Mux62;
output 	Mux621;
output 	Mux31;
output 	Mux32;
output 	Mux321;
output 	Mux0;
input 	Selector0;
input 	Mux241;
input 	Mux251;
input 	Mux261;
input 	Mux271;
input 	Mux410;
input 	Mux510;
input 	Mux64;
input 	Mux71;
input 	Mux291;
input 	Mux281;
input 	Mux301;
input 	Mux311;
input 	cuifRegSel_0;
input 	cuifRegSel_1;
input 	Selector68;
input 	Selector67;
input 	Selector64;
input 	Selector66;
input 	Selector65;
input 	Selector4;
input 	Selector41;
input 	Selector42;
input 	Selector1;
input 	Selector2;
input 	Selector3;
input 	Selector8;
input 	Selector9;
input 	Selector10;
input 	Selector11;
input 	Selector12;
input 	Selector13;
input 	Selector14;
input 	Selector15;
input 	Selector01;
input 	Mux231;
input 	Mux221;
input 	Mux211;
input 	Mux201;
input 	Mux191;
input 	Mux181;
input 	Mux171;
input 	Mux161;
input 	cuifRegSel_11;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \regs[21][0]~q ;
wire \regs[22][0]~q ;
wire \regs[26][1]~q ;
wire \regs[27][1]~q ;
wire \regs[1][1]~q ;
wire \regs[17][30]~q ;
wire \regs[18][30]~q ;
wire \regs[26][29]~q ;
wire \Mux37~2_combout ;
wire \regs[5][26]~q ;
wire \Mux5~10_combout ;
wire \regs[13][25]~q ;
wire \Mux6~17_combout ;
wire \regs[18][24]~q ;
wire \regs[24][24]~q ;
wire \Mux39~4_combout ;
wire \regs[5][24]~q ;
wire \Mux7~2_combout ;
wire \regs[16][23]~q ;
wire \regs[28][23]~q ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \regs[16][22]~q ;
wire \regs[5][22]~q ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux9~10_combout ;
wire \regs[18][21]~q ;
wire \Mux10~2_combout ;
wire \regs[8][19]~q ;
wire \regs[26][18]~q ;
wire \Mux45~4_combout ;
wire \regs[3][18]~q ;
wire \regs[13][18]~q ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \Mux13~10_combout ;
wire \Mux13~17_combout ;
wire \regs[8][17]~q ;
wire \regs[11][17]~q ;
wire \regs[17][15]~q ;
wire \regs[13][15]~q ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \Mux16~7_combout ;
wire \Mux16~17_combout ;
wire \regs[22][14]~q ;
wire \regs[26][14]~q ;
wire \Mux49~12_combout ;
wire \regs[13][14]~q ;
wire \Mux17~17_combout ;
wire \regs[3][13]~q ;
wire \regs[24][12]~q ;
wire \Mux19~0_combout ;
wire \regs[30][11]~q ;
wire \regs[13][11]~q ;
wire \Mux20~17_combout ;
wire \regs[22][10]~q ;
wire \regs[26][10]~q ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \regs[28][9]~q ;
wire \Mux22~10_combout ;
wire \regs[26][8]~q ;
wire \Mux55~2_combout ;
wire \regs[23][8]~q ;
wire \Mux56~2_combout ;
wire \regs[26][6]~q ;
wire \Mux57~2_combout ;
wire \regs[8][6]~q ;
wire \regs[17][5]~q ;
wire \regs[18][5]~q ;
wire \regs[30][5]~q ;
wire \regs[19][5]~q ;
wire \Mux26~0_combout ;
wire \Mux26~7_combout ;
wire \regs[24][4]~q ;
wire \regs[16][4]~q ;
wire \Mux59~4_combout ;
wire \Mux59~12_combout ;
wire \Mux27~4_combout ;
wire \Mux27~5_combout ;
wire \Mux27~14_combout ;
wire \Mux27~15_combout ;
wire \Mux60~4_combout ;
wire \regs[27][3]~q ;
wire \Mux28~14_combout ;
wire \Mux28~15_combout ;
wire \regs[4][31]~q ;
wire \regs[25][31]~q ;
wire \regs[27][31]~q ;
wire \regs~12_combout ;
wire \regs~15_combout ;
wire \regs~59_combout ;
wire \regs[21][0]~feeder_combout ;
wire \regs[26][1]~feeder_combout ;
wire \regs[27][1]~feeder_combout ;
wire \regs[18][30]~feeder_combout ;
wire \regs[17][30]~feeder_combout ;
wire \regs[26][29]~feeder_combout ;
wire \regs[5][24]~feeder_combout ;
wire \regs[8][19]~feeder_combout ;
wire \regs[11][17]~feeder_combout ;
wire \regs[8][17]~feeder_combout ;
wire \regs[17][15]~feeder_combout ;
wire \regs[22][14]~feeder_combout ;
wire \regs[26][14]~feeder_combout ;
wire \regs[3][13]~feeder_combout ;
wire \regs[24][12]~feeder_combout ;
wire \regs[30][11]~feeder_combout ;
wire \regs[22][10]~feeder_combout ;
wire \regs[26][10]~feeder_combout ;
wire \regs[28][9]~feeder_combout ;
wire \regs[23][8]~feeder_combout ;
wire \regs[8][6]~feeder_combout ;
wire \regs[19][5]~feeder_combout ;
wire \regs[18][5]~feeder_combout ;
wire \regs[30][5]~feeder_combout ;
wire \regs[27][3]~feeder_combout ;
wire \regs[25][31]~feeder_combout ;
wire \regs[27][31]~feeder_combout ;
wire \regs[4][31]~feeder_combout ;
wire \regs~4_combout ;
wire \regs~64_combout ;
wire \regs~5_combout ;
wire \regs[20][0]~feeder_combout ;
wire \Equal0~0_combout ;
wire \Decoder0~12_combout ;
wire \Decoder0~13_combout ;
wire \regs[20][0]~q ;
wire \Decoder0~16_combout ;
wire \regs[28][0]~q ;
wire \regs[24][0]~feeder_combout ;
wire \Decoder0~14_combout ;
wire \regs[24][0]~q ;
wire \Decoder0~15_combout ;
wire \regs[16][0]~q ;
wire \Mux63~4_combout ;
wire \Mux63~5_combout ;
wire \Decoder0~7_combout ;
wire \Decoder0~10_combout ;
wire \regs[18][0]~q ;
wire \Mux63~2_combout ;
wire \Decoder0~11_combout ;
wire \regs[30][0]~q ;
wire \Mux63~3_combout ;
wire \Mux63~6_combout ;
wire \Decoder0~0_combout ;
wire \Decoder0~1_combout ;
wire \Decoder0~2_combout ;
wire \regs[25][0]~q ;
wire \Decoder0~3_combout ;
wire \Decoder0~6_combout ;
wire \regs[29][0]~q ;
wire \regs[17][0]~feeder_combout ;
wire \Decoder0~5_combout ;
wire \regs[17][0]~q ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \Decoder0~17_combout ;
wire \Decoder0~18_combout ;
wire \regs[27][0]~q ;
wire \regs[31][0]~feeder_combout ;
wire \Decoder0~21_combout ;
wire \regs[31][0]~q ;
wire \regs[23][0]~feeder_combout ;
wire \Decoder0~19_combout ;
wire \regs[23][0]~q ;
wire \Mux63~7_combout ;
wire \Mux63~8_combout ;
wire \regs[9][0]~feeder_combout ;
wire \Decoder0~22_combout ;
wire \regs[9][0]~q ;
wire \Decoder0~25_combout ;
wire \Decoder0~26_combout ;
wire \regs[11][0]~q ;
wire \Decoder0~24_combout ;
wire \regs[8][0]~q ;
wire \Decoder0~23_combout ;
wire \regs[10][0]~q ;
wire \Mux63~10_combout ;
wire \Mux63~11_combout ;
wire \Decoder0~34_combout ;
wire \regs[14][0]~q ;
wire \Decoder0~37_combout ;
wire \regs[15][0]~q ;
wire \Decoder0~36_combout ;
wire \regs[12][0]~q ;
wire \Mux63~17_combout ;
wire \Mux63~18_combout ;
wire \Decoder0~29_combout ;
wire \regs[4][0]~q ;
wire \Decoder0~28_combout ;
wire \regs[5][0]~q ;
wire \Mux63~12_combout ;
wire \Decoder0~30_combout ;
wire \regs[7][0]~q ;
wire \Mux63~13_combout ;
wire \Decoder0~31_combout ;
wire \regs[1][0]~q ;
wire \Decoder0~33_combout ;
wire \regs[3][0]~q ;
wire \Mux63~14_combout ;
wire \Mux63~15_combout ;
wire \Mux63~16_combout ;
wire \Equal0~1_combout ;
wire \regs~6_combout ;
wire \regs~7_combout ;
wire \regs[31][1]~feeder_combout ;
wire \regs[31][1]~q ;
wire \regs[19][1]~feeder_combout ;
wire \Decoder0~20_combout ;
wire \regs[19][1]~q ;
wire \Mux30~7_combout ;
wire \Mux30~8_combout ;
wire \regs[29][1]~feeder_combout ;
wire \regs[29][1]~q ;
wire \regs[25][1]~feeder_combout ;
wire \regs[25][1]~q ;
wire \regs[21][1]~feeder_combout ;
wire \Decoder0~4_combout ;
wire \regs[21][1]~q ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \regs[18][1]~q ;
wire \Mux30~2_combout ;
wire \regs[22][1]~feeder_combout ;
wire \Decoder0~8_combout ;
wire \regs[22][1]~q ;
wire \Mux30~3_combout ;
wire \regs[28][1]~q ;
wire \regs[20][1]~q ;
wire \regs[24][1]~q ;
wire \Mux30~4_combout ;
wire \Mux30~5_combout ;
wire \Mux30~6_combout ;
wire \Mux30~9_combout ;
wire \regs[9][1]~q ;
wire \regs[10][1]~q ;
wire \Mux30~10_combout ;
wire \Mux30~11_combout ;
wire \regs[15][1]~q ;
wire \regs[14][1]~q ;
wire \regs[12][1]~q ;
wire \Decoder0~35_combout ;
wire \regs[13][1]~q ;
wire \Mux30~17_combout ;
wire \Mux30~18_combout ;
wire \regs[3][1]~q ;
wire \Mux30~14_combout ;
wire \Mux30~15_combout ;
wire \regs[7][1]~q ;
wire \Decoder0~27_combout ;
wire \regs[6][1]~q ;
wire \regs[5][1]~q ;
wire \Mux30~12_combout ;
wire \Mux30~13_combout ;
wire \Mux30~16_combout ;
wire \Mux30~19_combout ;
wire \regs~8_combout ;
wire \regs[31][30]~q ;
wire \regs[27][30]~q ;
wire \regs[23][30]~q ;
wire \Mux33~7_combout ;
wire \Mux33~8_combout ;
wire \regs[21][30]~q ;
wire \Mux33~0_combout ;
wire \regs[29][30]~q ;
wire \regs[25][30]~q ;
wire \Mux33~1_combout ;
wire \regs[16][30]~q ;
wire \regs[24][30]~q ;
wire \Mux33~4_combout ;
wire \regs[20][30]~q ;
wire \regs[28][30]~q ;
wire \Mux33~5_combout ;
wire \regs[22][30]~feeder_combout ;
wire \regs[22][30]~q ;
wire \Decoder0~9_combout ;
wire \regs[26][30]~q ;
wire \Mux33~2_combout ;
wire \Mux33~3_combout ;
wire \Mux33~6_combout ;
wire \regs[14][30]~q ;
wire \regs[15][30]~q ;
wire \regs[13][30]~q ;
wire \regs[12][30]~q ;
wire \Mux33~17_combout ;
wire \Mux33~18_combout ;
wire \regs[10][30]~q ;
wire \Mux33~10_combout ;
wire \regs[11][30]~feeder_combout ;
wire \regs[11][30]~q ;
wire \regs[9][30]~q ;
wire \Mux33~11_combout ;
wire \regs[6][30]~q ;
wire \regs[7][30]~q ;
wire \regs[4][30]~q ;
wire \Mux33~12_combout ;
wire \Mux33~13_combout ;
wire \Decoder0~32_combout ;
wire \regs[2][30]~q ;
wire \regs[3][30]~feeder_combout ;
wire \regs[3][30]~q ;
wire \regs[1][30]~q ;
wire \Mux33~14_combout ;
wire \Mux33~15_combout ;
wire \Mux33~16_combout ;
wire \Mux1~14_combout ;
wire \Mux1~15_combout ;
wire \regs[8][30]~feeder_combout ;
wire \regs[8][30]~q ;
wire \Mux1~12_combout ;
wire \Mux1~13_combout ;
wire \Mux1~16_combout ;
wire \Mux1~17_combout ;
wire \Mux1~18_combout ;
wire \regs[5][30]~q ;
wire \Mux1~10_combout ;
wire \Mux1~11_combout ;
wire \Mux1~19_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \regs[19][30]~q ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \regs[30][30]~feeder_combout ;
wire \regs[30][30]~q ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \Mux1~9_combout ;
wire \regs~9_combout ;
wire \regs[31][29]~q ;
wire \regs[23][29]~feeder_combout ;
wire \regs[23][29]~q ;
wire \regs[27][29]~feeder_combout ;
wire \regs[27][29]~q ;
wire \Mux34~7_combout ;
wire \Mux34~8_combout ;
wire \regs[21][29]~feeder_combout ;
wire \regs[21][29]~q ;
wire \regs[25][29]~q ;
wire \Mux34~0_combout ;
wire \regs[29][29]~q ;
wire \Mux34~1_combout ;
wire \regs[28][29]~q ;
wire \regs[24][29]~q ;
wire \regs[20][29]~q ;
wire \Mux34~4_combout ;
wire \Mux34~5_combout ;
wire \regs[30][29]~q ;
wire \regs[22][29]~q ;
wire \Mux34~2_combout ;
wire \Mux34~3_combout ;
wire \Mux34~6_combout ;
wire \regs[5][29]~q ;
wire \Mux34~10_combout ;
wire \regs[7][29]~q ;
wire \regs[6][29]~q ;
wire \Mux34~11_combout ;
wire \regs[14][29]~q ;
wire \regs[13][29]~q ;
wire \regs[12][29]~q ;
wire \Mux34~17_combout ;
wire \regs[15][29]~q ;
wire \Mux34~18_combout ;
wire \regs[3][29]~q ;
wire \regs[1][29]~q ;
wire \Mux34~14_combout ;
wire \regs[2][29]~q ;
wire \Mux34~15_combout ;
wire \regs[9][29]~q ;
wire \regs[11][29]~q ;
wire \regs[8][29]~q ;
wire \Mux34~12_combout ;
wire \Mux34~13_combout ;
wire \Mux34~16_combout ;
wire \regs[16][29]~q ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \regs[18][29]~q ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \Mux2~6_combout ;
wire \regs[19][29]~q ;
wire \Mux2~7_combout ;
wire \Mux2~8_combout ;
wire \regs[17][29]~q ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~9_combout ;
wire \Mux2~17_combout ;
wire \Mux2~18_combout ;
wire \regs[10][29]~q ;
wire \Mux2~10_combout ;
wire \Mux2~11_combout ;
wire \Mux2~14_combout ;
wire \Mux2~15_combout ;
wire \regs[4][29]~q ;
wire \Mux2~12_combout ;
wire \Mux2~13_combout ;
wire \Mux2~16_combout ;
wire \Mux2~19_combout ;
wire \regs~10_combout ;
wire \regs[30][28]~q ;
wire \regs[18][28]~q ;
wire \Mux35~2_combout ;
wire \Mux35~3_combout ;
wire \regs[20][28]~q ;
wire \regs[28][28]~q ;
wire \regs[24][28]~q ;
wire \regs[16][28]~q ;
wire \Mux35~4_combout ;
wire \Mux35~5_combout ;
wire \Mux35~6_combout ;
wire \regs[27][28]~q ;
wire \regs[31][28]~feeder_combout ;
wire \regs[31][28]~q ;
wire \regs[19][28]~feeder_combout ;
wire \regs[19][28]~q ;
wire \Mux35~7_combout ;
wire \Mux35~8_combout ;
wire \regs[29][28]~feeder_combout ;
wire \regs[29][28]~q ;
wire \regs[25][28]~q ;
wire \regs[17][28]~feeder_combout ;
wire \regs[17][28]~q ;
wire \Mux35~0_combout ;
wire \Mux35~1_combout ;
wire \regs[14][28]~q ;
wire \regs[13][28]~feeder_combout ;
wire \regs[13][28]~q ;
wire \regs[12][28]~q ;
wire \Mux35~17_combout ;
wire \regs[15][28]~q ;
wire \Mux35~18_combout ;
wire \regs[9][28]~q ;
wire \regs[11][28]~q ;
wire \regs[10][28]~q ;
wire \regs[8][28]~q ;
wire \Mux35~10_combout ;
wire \Mux35~11_combout ;
wire \regs[2][28]~q ;
wire \regs[1][28]~q ;
wire \Mux35~14_combout ;
wire \Mux35~15_combout ;
wire \regs[6][28]~q ;
wire \regs[7][28]~q ;
wire \regs[4][28]~q ;
wire \Mux35~12_combout ;
wire \Mux35~13_combout ;
wire \Mux35~16_combout ;
wire \Mux3~17_combout ;
wire \Mux3~18_combout ;
wire \Mux3~12_combout ;
wire \Mux3~13_combout ;
wire \regs[3][28]~feeder_combout ;
wire \regs[3][28]~q ;
wire \Mux3~14_combout ;
wire \Mux3~15_combout ;
wire \Mux3~16_combout ;
wire \regs[5][28]~q ;
wire \Mux3~10_combout ;
wire \Mux3~11_combout ;
wire \Mux3~19_combout ;
wire \regs[23][28]~feeder_combout ;
wire \regs[23][28]~q ;
wire \Mux3~7_combout ;
wire \Mux3~8_combout ;
wire \regs[21][28]~feeder_combout ;
wire \regs[21][28]~q ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \regs[26][28]~feeder_combout ;
wire \regs[26][28]~q ;
wire \regs[22][28]~q ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \Mux3~6_combout ;
wire \Mux3~9_combout ;
wire \regs~11_combout ;
wire \regs~13_combout ;
wire \regs[20][27]~feeder_combout ;
wire \regs[20][27]~q ;
wire \regs[16][27]~q ;
wire \Mux36~4_combout ;
wire \regs[28][27]~q ;
wire \Mux36~5_combout ;
wire \regs[30][27]~q ;
wire \regs[18][27]~q ;
wire \Mux36~2_combout ;
wire \Mux36~3_combout ;
wire \Mux36~6_combout ;
wire \regs[23][27]~feeder_combout ;
wire \regs[23][27]~q ;
wire \regs[31][27]~feeder_combout ;
wire \regs[31][27]~q ;
wire \regs[27][27]~q ;
wire \Mux36~7_combout ;
wire \Mux36~8_combout ;
wire \regs[21][27]~feeder_combout ;
wire \regs[21][27]~q ;
wire \regs[29][27]~q ;
wire \regs[25][27]~q ;
wire \regs[17][27]~q ;
wire \Mux36~0_combout ;
wire \Mux36~1_combout ;
wire \regs[6][27]~q ;
wire \regs[7][27]~q ;
wire \regs[4][27]~q ;
wire \Mux36~10_combout ;
wire \Mux36~11_combout ;
wire \regs[2][27]~q ;
wire \regs[3][27]~q ;
wire \regs[1][27]~q ;
wire \Mux36~14_combout ;
wire \Mux36~15_combout ;
wire \regs[8][27]~q ;
wire \regs[10][27]~feeder_combout ;
wire \regs[10][27]~q ;
wire \Mux36~12_combout ;
wire \regs[11][27]~q ;
wire \regs[9][27]~q ;
wire \Mux36~13_combout ;
wire \Mux36~16_combout ;
wire \regs[14][27]~q ;
wire \regs[15][27]~q ;
wire \regs[13][27]~q ;
wire \regs[12][27]~q ;
wire \Mux36~17_combout ;
wire \Mux36~18_combout ;
wire \regs[19][27]~feeder_combout ;
wire \regs[19][27]~q ;
wire \Mux4~7_combout ;
wire \Mux4~8_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \regs[22][27]~feeder_combout ;
wire \regs[22][27]~q ;
wire \regs[26][27]~q ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \regs[24][27]~q ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Mux4~6_combout ;
wire \Mux4~9_combout ;
wire \Mux4~17_combout ;
wire \Mux4~18_combout ;
wire \Mux4~10_combout ;
wire \Mux4~11_combout ;
wire \Mux4~14_combout ;
wire \Mux4~15_combout ;
wire \regs[5][27]~q ;
wire \Mux4~12_combout ;
wire \Mux4~13_combout ;
wire \Mux4~16_combout ;
wire \Mux4~19_combout ;
wire \regs~14_combout ;
wire \regs~16_combout ;
wire \regs[20][26]~q ;
wire \regs[28][26]~q ;
wire \regs[24][26]~q ;
wire \regs[16][26]~q ;
wire \Mux37~4_combout ;
wire \Mux37~5_combout ;
wire \regs[30][26]~q ;
wire \regs[22][26]~q ;
wire \Mux37~3_combout ;
wire \Mux37~6_combout ;
wire \regs[27][26]~feeder_combout ;
wire \regs[27][26]~q ;
wire \regs[31][26]~q ;
wire \regs[23][26]~q ;
wire \regs[19][26]~q ;
wire \Mux37~7_combout ;
wire \Mux37~8_combout ;
wire \regs[25][26]~q ;
wire \regs[29][26]~q ;
wire \regs[21][26]~feeder_combout ;
wire \regs[21][26]~q ;
wire \regs[17][26]~q ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \regs[9][26]~q ;
wire \regs[11][26]~q ;
wire \regs[10][26]~q ;
wire \regs[8][26]~q ;
wire \Mux37~10_combout ;
wire \Mux37~11_combout ;
wire \regs[14][26]~q ;
wire \regs[15][26]~q ;
wire \regs[12][26]~q ;
wire \Mux37~17_combout ;
wire \Mux37~18_combout ;
wire \regs[6][26]~q ;
wire \regs[7][26]~q ;
wire \regs[4][26]~q ;
wire \Mux37~12_combout ;
wire \Mux37~13_combout ;
wire \regs[2][26]~q ;
wire \regs[3][26]~q ;
wire \regs[1][26]~q ;
wire \Mux37~14_combout ;
wire \Mux37~15_combout ;
wire \Mux37~16_combout ;
wire \Mux5~7_combout ;
wire \Mux5~8_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \regs[26][26]~q ;
wire \regs[18][26]~q ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux5~4_combout ;
wire \Mux5~5_combout ;
wire \Mux5~6_combout ;
wire \Mux5~9_combout ;
wire \Mux5~12_combout ;
wire \Mux5~13_combout ;
wire \Mux5~14_combout ;
wire \Mux5~15_combout ;
wire \Mux5~16_combout ;
wire \regs[13][26]~q ;
wire \Mux5~17_combout ;
wire \Mux5~18_combout ;
wire \Mux5~11_combout ;
wire \Mux5~19_combout ;
wire \regs~17_combout ;
wire \regs~18_combout ;
wire \regs~19_combout ;
wire \regs[28][25]~q ;
wire \regs[20][25]~q ;
wire \regs[16][25]~q ;
wire \Mux38~4_combout ;
wire \Mux38~5_combout ;
wire \regs[30][25]~q ;
wire \regs[18][25]~q ;
wire \Mux38~2_combout ;
wire \Mux38~3_combout ;
wire \Mux38~6_combout ;
wire \regs[21][25]~feeder_combout ;
wire \regs[21][25]~q ;
wire \regs[25][25]~q ;
wire \regs[17][25]~q ;
wire \Mux38~0_combout ;
wire \regs[29][25]~q ;
wire \Mux38~1_combout ;
wire \regs[31][25]~feeder_combout ;
wire \regs[31][25]~q ;
wire \regs[23][25]~q ;
wire \regs[27][25]~feeder_combout ;
wire \regs[27][25]~q ;
wire \Mux38~7_combout ;
wire \Mux38~8_combout ;
wire \regs[6][25]~q ;
wire \regs[4][25]~q ;
wire \Mux38~10_combout ;
wire \regs[7][25]~q ;
wire \Mux38~11_combout ;
wire \regs[14][25]~q ;
wire \regs[15][25]~q ;
wire \regs[12][25]~q ;
wire \Mux38~17_combout ;
wire \Mux38~18_combout ;
wire \regs[9][25]~q ;
wire \regs[11][25]~q ;
wire \regs[8][25]~q ;
wire \Mux38~12_combout ;
wire \Mux38~13_combout ;
wire \regs[3][25]~feeder_combout ;
wire \regs[3][25]~q ;
wire \regs[1][25]~q ;
wire \Mux38~14_combout ;
wire \regs[2][25]~q ;
wire \Mux38~15_combout ;
wire \Mux38~16_combout ;
wire \regs[24][25]~q ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \regs[22][25]~feeder_combout ;
wire \regs[22][25]~q ;
wire \regs[26][25]~q ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \Mux6~6_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \regs[19][25]~feeder_combout ;
wire \regs[19][25]~q ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \Mux6~9_combout ;
wire \Mux6~18_combout ;
wire \regs[10][25]~q ;
wire \Mux6~10_combout ;
wire \Mux6~11_combout ;
wire \Mux6~14_combout ;
wire \Mux6~15_combout ;
wire \regs[5][25]~q ;
wire \Mux6~12_combout ;
wire \Mux6~13_combout ;
wire \Mux6~16_combout ;
wire \Mux6~19_combout ;
wire \regs~20_combout ;
wire \regs~21_combout ;
wire \regs~22_combout ;
wire \regs[31][24]~q ;
wire \regs[27][24]~q ;
wire \regs[19][24]~q ;
wire \regs[23][24]~q ;
wire \Mux39~7_combout ;
wire \Mux39~8_combout ;
wire \regs[29][24]~q ;
wire \regs[25][24]~q ;
wire \regs[21][24]~q ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \regs[28][24]~q ;
wire \regs[20][24]~q ;
wire \Mux39~5_combout ;
wire \regs[22][24]~q ;
wire \regs[26][24]~q ;
wire \Mux39~2_combout ;
wire \Mux39~3_combout ;
wire \Mux39~6_combout ;
wire \regs[14][24]~feeder_combout ;
wire \regs[14][24]~q ;
wire \regs[15][24]~q ;
wire \regs[12][24]~q ;
wire \Mux39~17_combout ;
wire \Mux39~18_combout ;
wire \regs[10][24]~q ;
wire \Mux39~10_combout ;
wire \regs[11][24]~q ;
wire \regs[9][24]~q ;
wire \Mux39~11_combout ;
wire \regs[3][24]~q ;
wire \regs[1][24]~q ;
wire \Mux39~14_combout ;
wire \regs[2][24]~q ;
wire \Mux39~15_combout ;
wire \regs[4][24]~q ;
wire \Mux39~12_combout ;
wire \regs[7][24]~q ;
wire \Mux39~13_combout ;
wire \Mux39~16_combout ;
wire \regs[30][24]~q ;
wire \Mux7~3_combout ;
wire \regs[16][24]~q ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \Mux7~6_combout ;
wire \regs[17][24]~q ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux7~7_combout ;
wire \Mux7~8_combout ;
wire \Mux7~9_combout ;
wire \regs[6][24]~feeder_combout ;
wire \regs[6][24]~q ;
wire \Mux7~10_combout ;
wire \Mux7~11_combout ;
wire \regs[13][24]~feeder_combout ;
wire \regs[13][24]~q ;
wire \Mux7~17_combout ;
wire \Mux7~18_combout ;
wire \regs[8][24]~q ;
wire \Mux7~12_combout ;
wire \Mux7~13_combout ;
wire \Mux7~14_combout ;
wire \Mux7~15_combout ;
wire \Mux7~16_combout ;
wire \Mux7~19_combout ;
wire \regs~23_combout ;
wire \regs[29][23]~q ;
wire \regs[21][23]~feeder_combout ;
wire \regs[21][23]~q ;
wire \regs[25][23]~feeder_combout ;
wire \regs[25][23]~q ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \regs[26][23]~q ;
wire \regs[18][23]~q ;
wire \Mux40~2_combout ;
wire \Mux40~3_combout ;
wire \regs[24][23]~q ;
wire \regs[20][23]~q ;
wire \Mux40~4_combout ;
wire \Mux40~5_combout ;
wire \Mux40~6_combout ;
wire \regs[31][23]~q ;
wire \regs[23][23]~feeder_combout ;
wire \regs[23][23]~q ;
wire \regs[27][23]~feeder_combout ;
wire \regs[27][23]~q ;
wire \Mux40~7_combout ;
wire \Mux40~8_combout ;
wire \regs[7][23]~q ;
wire \regs[6][23]~q ;
wire \regs[5][23]~q ;
wire \Mux40~10_combout ;
wire \Mux40~11_combout ;
wire \regs[14][23]~feeder_combout ;
wire \regs[14][23]~q ;
wire \regs[15][23]~q ;
wire \regs[12][23]~q ;
wire \Mux40~17_combout ;
wire \Mux40~18_combout ;
wire \regs[2][23]~q ;
wire \regs[1][23]~q ;
wire \Mux40~14_combout ;
wire \Mux40~15_combout ;
wire \regs[8][23]~q ;
wire \Mux40~12_combout ;
wire \regs[11][23]~q ;
wire \regs[9][23]~q ;
wire \Mux40~13_combout ;
wire \Mux40~16_combout ;
wire \regs[22][23]~feeder_combout ;
wire \regs[22][23]~q ;
wire \regs[30][23]~q ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Mux8~6_combout ;
wire \regs[19][23]~q ;
wire \Mux8~7_combout ;
wire \Mux8~8_combout ;
wire \regs[17][23]~q ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux8~9_combout ;
wire \regs[13][23]~feeder_combout ;
wire \regs[13][23]~q ;
wire \Mux8~17_combout ;
wire \Mux8~18_combout ;
wire \regs[10][23]~q ;
wire \Mux8~10_combout ;
wire \Mux8~11_combout ;
wire \regs[3][23]~feeder_combout ;
wire \regs[3][23]~q ;
wire \Mux8~14_combout ;
wire \Mux8~15_combout ;
wire \regs[4][23]~q ;
wire \Mux8~12_combout ;
wire \Mux8~13_combout ;
wire \Mux8~16_combout ;
wire \Mux8~19_combout ;
wire \regs~24_combout ;
wire \regs[29][22]~feeder_combout ;
wire \regs[29][22]~q ;
wire \regs[25][22]~q ;
wire \regs[21][22]~q ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \regs[27][22]~feeder_combout ;
wire \regs[27][22]~q ;
wire \regs[31][22]~q ;
wire \regs[23][22]~feeder_combout ;
wire \regs[23][22]~q ;
wire \Mux41~7_combout ;
wire \Mux41~8_combout ;
wire \regs[28][22]~q ;
wire \regs[20][22]~q ;
wire \regs[24][22]~q ;
wire \Mux41~4_combout ;
wire \Mux41~5_combout ;
wire \regs[22][22]~feeder_combout ;
wire \regs[22][22]~q ;
wire \regs[26][22]~q ;
wire \Mux41~2_combout ;
wire \Mux41~3_combout ;
wire \Mux41~6_combout ;
wire \regs[11][22]~q ;
wire \regs[9][22]~q ;
wire \regs[10][22]~q ;
wire \Mux41~10_combout ;
wire \Mux41~11_combout ;
wire \regs[7][22]~q ;
wire \regs[4][22]~q ;
wire \Mux41~12_combout ;
wire \Mux41~13_combout ;
wire \regs[2][22]~q ;
wire \regs[1][22]~q ;
wire \Mux41~14_combout ;
wire \Mux41~15_combout ;
wire \Mux41~16_combout ;
wire \regs[14][22]~feeder_combout ;
wire \regs[14][22]~q ;
wire \regs[15][22]~feeder_combout ;
wire \regs[15][22]~q ;
wire \regs[12][22]~q ;
wire \Mux41~17_combout ;
wire \Mux41~18_combout ;
wire \regs[30][22]~q ;
wire \regs[18][22]~q ;
wire \Mux9~2_combout ;
wire \Mux9~3_combout ;
wire \Mux9~6_combout ;
wire \regs[17][22]~q ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \regs[19][22]~q ;
wire \Mux9~7_combout ;
wire \Mux9~8_combout ;
wire \Mux9~9_combout ;
wire \regs[6][22]~q ;
wire \Mux9~11_combout ;
wire \regs[13][22]~q ;
wire \Mux9~17_combout ;
wire \Mux9~18_combout ;
wire \regs[3][22]~feeder_combout ;
wire \regs[3][22]~q ;
wire \Mux9~14_combout ;
wire \Mux9~15_combout ;
wire \regs[8][22]~q ;
wire \Mux9~12_combout ;
wire \Mux9~13_combout ;
wire \Mux9~16_combout ;
wire \Mux9~19_combout ;
wire \regs~25_combout ;
wire \regs[23][21]~feeder_combout ;
wire \regs[23][21]~q ;
wire \regs[31][21]~q ;
wire \regs[27][21]~feeder_combout ;
wire \regs[27][21]~q ;
wire \Mux42~7_combout ;
wire \Mux42~8_combout ;
wire \regs[21][21]~feeder_combout ;
wire \regs[21][21]~q ;
wire \regs[29][21]~feeder_combout ;
wire \regs[29][21]~q ;
wire \regs[17][21]~feeder_combout ;
wire \regs[17][21]~q ;
wire \regs[25][21]~feeder_combout ;
wire \regs[25][21]~q ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \regs[24][21]~q ;
wire \regs[20][21]~q ;
wire \Mux42~4_combout ;
wire \Mux42~5_combout ;
wire \regs[26][21]~q ;
wire \regs[22][21]~q ;
wire \Mux42~2_combout ;
wire \Mux42~3_combout ;
wire \Mux42~6_combout ;
wire \regs[3][21]~feeder_combout ;
wire \regs[3][21]~q ;
wire \regs[1][21]~q ;
wire \Mux42~14_combout ;
wire \regs[2][21]~q ;
wire \Mux42~15_combout ;
wire \regs[9][21]~feeder_combout ;
wire \regs[9][21]~q ;
wire \regs[11][21]~q ;
wire \regs[8][21]~feeder_combout ;
wire \regs[8][21]~q ;
wire \Mux42~12_combout ;
wire \Mux42~13_combout ;
wire \Mux42~16_combout ;
wire \regs[5][21]~q ;
wire \Mux42~10_combout ;
wire \regs[7][21]~q ;
wire \regs[6][21]~q ;
wire \Mux42~11_combout ;
wire \regs[12][21]~q ;
wire \Mux42~17_combout ;
wire \regs[14][21]~q ;
wire \regs[15][21]~q ;
wire \Mux42~18_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \regs[28][21]~q ;
wire \regs[16][21]~q ;
wire \Mux10~4_combout ;
wire \Mux10~5_combout ;
wire \regs[30][21]~q ;
wire \Mux10~3_combout ;
wire \Mux10~6_combout ;
wire \regs[19][21]~q ;
wire \Mux10~7_combout ;
wire \Mux10~8_combout ;
wire \Mux10~9_combout ;
wire \regs[13][21]~q ;
wire \Mux10~17_combout ;
wire \Mux10~18_combout ;
wire \regs[10][21]~q ;
wire \Mux10~10_combout ;
wire \Mux10~11_combout ;
wire \Mux10~14_combout ;
wire \Mux10~15_combout ;
wire \regs[4][21]~q ;
wire \Mux10~12_combout ;
wire \Mux10~13_combout ;
wire \Mux10~16_combout ;
wire \Mux10~19_combout ;
wire \regs~26_combout ;
wire \regs[27][20]~feeder_combout ;
wire \regs[27][20]~q ;
wire \regs[31][20]~q ;
wire \regs[23][20]~q ;
wire \regs[19][20]~q ;
wire \Mux43~7_combout ;
wire \Mux43~8_combout ;
wire \regs[28][20]~q ;
wire \regs[16][20]~q ;
wire \Mux43~4_combout ;
wire \Mux43~5_combout ;
wire \regs[30][20]~q ;
wire \regs[18][20]~q ;
wire \Mux43~2_combout ;
wire \Mux43~3_combout ;
wire \Mux43~6_combout ;
wire \regs[25][20]~q ;
wire \regs[29][20]~feeder_combout ;
wire \regs[29][20]~q ;
wire \regs[21][20]~feeder_combout ;
wire \regs[21][20]~q ;
wire \regs[17][20]~q ;
wire \Mux43~0_combout ;
wire \Mux43~1_combout ;
wire \regs[14][20]~feeder_combout ;
wire \regs[14][20]~q ;
wire \regs[15][20]~q ;
wire \regs[12][20]~q ;
wire \Mux43~17_combout ;
wire \Mux43~18_combout ;
wire \regs[9][20]~feeder_combout ;
wire \regs[9][20]~q ;
wire \regs[11][20]~q ;
wire \regs[8][20]~feeder_combout ;
wire \regs[8][20]~q ;
wire \regs[10][20]~q ;
wire \Mux43~10_combout ;
wire \Mux43~11_combout ;
wire \regs[2][20]~q ;
wire \regs[1][20]~q ;
wire \Mux43~14_combout ;
wire \Mux43~15_combout ;
wire \regs[6][20]~feeder_combout ;
wire \regs[6][20]~q ;
wire \regs[7][20]~q ;
wire \regs[5][20]~feeder_combout ;
wire \regs[5][20]~q ;
wire \regs[4][20]~q ;
wire \Mux43~12_combout ;
wire \Mux43~13_combout ;
wire \Mux43~16_combout ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \regs[24][20]~feeder_combout ;
wire \regs[24][20]~q ;
wire \regs[20][20]~q ;
wire \Mux11~4_combout ;
wire \Mux11~5_combout ;
wire \regs[26][20]~q ;
wire \regs[22][20]~q ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \Mux11~6_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux11~9_combout ;
wire \Mux11~10_combout ;
wire \Mux11~11_combout ;
wire \regs[13][20]~feeder_combout ;
wire \regs[13][20]~q ;
wire \Mux11~17_combout ;
wire \Mux11~18_combout ;
wire \regs[3][20]~q ;
wire \Mux11~14_combout ;
wire \Mux11~15_combout ;
wire \Mux11~12_combout ;
wire \Mux11~13_combout ;
wire \Mux11~16_combout ;
wire \Mux11~19_combout ;
wire \regs~27_combout ;
wire \regs[23][19]~q ;
wire \regs[31][19]~q ;
wire \regs[27][19]~feeder_combout ;
wire \regs[27][19]~q ;
wire \Mux44~7_combout ;
wire \Mux44~8_combout ;
wire \regs[24][19]~feeder_combout ;
wire \regs[24][19]~q ;
wire \regs[28][19]~q ;
wire \regs[16][19]~q ;
wire \Mux44~4_combout ;
wire \Mux44~5_combout ;
wire \regs[26][19]~q ;
wire \regs[30][19]~q ;
wire \regs[18][19]~q ;
wire \Mux44~2_combout ;
wire \Mux44~3_combout ;
wire \Mux44~6_combout ;
wire \regs[29][19]~feeder_combout ;
wire \regs[29][19]~q ;
wire \regs[21][19]~q ;
wire \regs[25][19]~feeder_combout ;
wire \regs[25][19]~q ;
wire \regs[17][19]~q ;
wire \Mux44~0_combout ;
wire \Mux44~1_combout ;
wire \regs[14][19]~q ;
wire \regs[15][19]~q ;
wire \regs[13][19]~q ;
wire \Mux44~17_combout ;
wire \Mux44~18_combout ;
wire \regs[2][19]~q ;
wire \regs[3][19]~q ;
wire \regs[1][19]~q ;
wire \Mux44~14_combout ;
wire \Mux44~15_combout ;
wire \regs[9][19]~feeder_combout ;
wire \regs[9][19]~q ;
wire \regs[11][19]~q ;
wire \regs[10][19]~q ;
wire \Mux44~12_combout ;
wire \Mux44~13_combout ;
wire \Mux44~16_combout ;
wire \regs[6][19]~q ;
wire \regs[7][19]~feeder_combout ;
wire \regs[7][19]~q ;
wire \regs[5][19]~q ;
wire \Mux44~10_combout ;
wire \Mux44~11_combout ;
wire \regs[20][19]~q ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \regs[22][19]~feeder_combout ;
wire \regs[22][19]~q ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Mux12~6_combout ;
wire \regs[19][19]~feeder_combout ;
wire \regs[19][19]~q ;
wire \Mux12~7_combout ;
wire \Mux12~8_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux12~9_combout ;
wire \Mux12~10_combout ;
wire \Mux12~11_combout ;
wire \regs[12][19]~feeder_combout ;
wire \regs[12][19]~q ;
wire \Mux12~17_combout ;
wire \Mux12~18_combout ;
wire \regs[4][19]~q ;
wire \Mux12~12_combout ;
wire \Mux12~13_combout ;
wire \Mux12~14_combout ;
wire \Mux12~15_combout ;
wire \Mux12~16_combout ;
wire \Mux12~19_combout ;
wire \regs~28_combout ;
wire \regs[22][18]~feeder_combout ;
wire \regs[22][18]~q ;
wire \regs[30][18]~q ;
wire \regs[18][18]~q ;
wire \Mux45~2_combout ;
wire \Mux45~3_combout ;
wire \regs[20][18]~q ;
wire \regs[28][18]~q ;
wire \Mux45~5_combout ;
wire \Mux45~6_combout ;
wire \regs[27][18]~q ;
wire \regs[31][18]~q ;
wire \regs[23][18]~q ;
wire \regs[19][18]~q ;
wire \Mux45~7_combout ;
wire \Mux45~8_combout ;
wire \regs[25][18]~q ;
wire \regs[29][18]~q ;
wire \regs[21][18]~q ;
wire \regs[17][18]~q ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \regs[14][18]~q ;
wire \regs[15][18]~q ;
wire \regs[12][18]~q ;
wire \Mux45~17_combout ;
wire \Mux45~18_combout ;
wire \regs[9][18]~q ;
wire \regs[11][18]~q ;
wire \regs[8][18]~q ;
wire \Mux45~10_combout ;
wire \Mux45~11_combout ;
wire \regs[2][18]~q ;
wire \regs[1][18]~q ;
wire \Mux45~14_combout ;
wire \Mux45~15_combout ;
wire \regs[7][18]~q ;
wire \regs[5][18]~feeder_combout ;
wire \regs[5][18]~q ;
wire \regs[4][18]~q ;
wire \Mux45~12_combout ;
wire \Mux45~13_combout ;
wire \Mux45~16_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux13~7_combout ;
wire \Mux13~8_combout ;
wire \regs[24][18]~q ;
wire \regs[16][18]~q ;
wire \Mux13~4_combout ;
wire \Mux13~5_combout ;
wire \Mux13~6_combout ;
wire \Mux13~9_combout ;
wire \regs[6][18]~feeder_combout ;
wire \regs[6][18]~q ;
wire \Mux13~11_combout ;
wire \Mux13~18_combout ;
wire \Mux13~14_combout ;
wire \Mux13~15_combout ;
wire \regs[10][18]~q ;
wire \Mux13~12_combout ;
wire \Mux13~13_combout ;
wire \Mux13~16_combout ;
wire \Mux13~19_combout ;
wire \regs~29_combout ;
wire \regs[21][17]~q ;
wire \regs[29][17]~q ;
wire \regs[17][17]~feeder_combout ;
wire \regs[17][17]~q ;
wire \Mux46~0_combout ;
wire \Mux46~1_combout ;
wire \regs[23][17]~q ;
wire \regs[31][17]~q ;
wire \regs[19][17]~q ;
wire \Mux46~7_combout ;
wire \Mux46~8_combout ;
wire \regs[16][17]~q ;
wire \Mux46~4_combout ;
wire \regs[28][17]~q ;
wire \Mux46~5_combout ;
wire \regs[30][17]~q ;
wire \regs[18][17]~q ;
wire \Mux46~2_combout ;
wire \Mux46~3_combout ;
wire \Mux46~6_combout ;
wire \regs[14][17]~q ;
wire \regs[15][17]~q ;
wire \regs[12][17]~q ;
wire \Mux46~17_combout ;
wire \Mux46~18_combout ;
wire \regs[4][17]~feeder_combout ;
wire \regs[4][17]~q ;
wire \Mux46~10_combout ;
wire \regs[6][17]~q ;
wire \regs[7][17]~q ;
wire \Mux46~11_combout ;
wire \regs[9][17]~feeder_combout ;
wire \regs[9][17]~q ;
wire \regs[10][17]~q ;
wire \Mux46~12_combout ;
wire \Mux46~13_combout ;
wire \regs[2][17]~feeder_combout ;
wire \regs[2][17]~q ;
wire \regs[3][17]~q ;
wire \regs[1][17]~q ;
wire \Mux46~14_combout ;
wire \Mux46~15_combout ;
wire \Mux46~16_combout ;
wire \regs[27][17]~q ;
wire \Mux14~7_combout ;
wire \Mux14~8_combout ;
wire \regs[20][17]~q ;
wire \regs[24][17]~q ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \regs[22][17]~q ;
wire \regs[26][17]~feeder_combout ;
wire \regs[26][17]~q ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \Mux14~6_combout ;
wire \regs[25][17]~q ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Mux14~9_combout ;
wire \Mux14~10_combout ;
wire \Mux14~11_combout ;
wire \regs[13][17]~q ;
wire \Mux14~17_combout ;
wire \Mux14~18_combout ;
wire \Mux14~14_combout ;
wire \Mux14~15_combout ;
wire \regs[5][17]~q ;
wire \Mux14~12_combout ;
wire \Mux14~13_combout ;
wire \Mux14~16_combout ;
wire \Mux14~19_combout ;
wire \regs~30_combout ;
wire \regs[25][16]~q ;
wire \regs[29][16]~q ;
wire \regs[21][16]~feeder_combout ;
wire \regs[21][16]~q ;
wire \regs[17][16]~q ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \regs[22][16]~feeder_combout ;
wire \regs[22][16]~q ;
wire \regs[30][16]~q ;
wire \regs[18][16]~q ;
wire \Mux47~2_combout ;
wire \Mux47~3_combout ;
wire \regs[20][16]~q ;
wire \regs[28][16]~q ;
wire \regs[24][16]~feeder_combout ;
wire \regs[24][16]~q ;
wire \regs[16][16]~q ;
wire \Mux47~4_combout ;
wire \Mux47~5_combout ;
wire \Mux47~6_combout ;
wire \regs[27][16]~feeder_combout ;
wire \regs[27][16]~q ;
wire \regs[31][16]~q ;
wire \regs[23][16]~q ;
wire \regs[19][16]~q ;
wire \Mux47~7_combout ;
wire \Mux47~8_combout ;
wire \regs[14][16]~q ;
wire \regs[15][16]~feeder_combout ;
wire \regs[15][16]~q ;
wire \regs[12][16]~q ;
wire \Mux47~17_combout ;
wire \Mux47~18_combout ;
wire \regs[9][16]~feeder_combout ;
wire \regs[9][16]~q ;
wire \regs[11][16]~q ;
wire \regs[10][16]~q ;
wire \regs[8][16]~q ;
wire \Mux47~10_combout ;
wire \Mux47~11_combout ;
wire \regs[2][16]~q ;
wire \regs[1][16]~q ;
wire \Mux47~14_combout ;
wire \Mux47~15_combout ;
wire \regs[6][16]~q ;
wire \regs[7][16]~q ;
wire \regs[5][16]~q ;
wire \regs[4][16]~q ;
wire \Mux47~12_combout ;
wire \Mux47~13_combout ;
wire \Mux47~16_combout ;
wire \regs[13][16]~q ;
wire \Mux15~17_combout ;
wire \Mux15~18_combout ;
wire \Mux15~10_combout ;
wire \Mux15~11_combout ;
wire \regs[3][16]~q ;
wire \Mux15~14_combout ;
wire \Mux15~15_combout ;
wire \Mux15~12_combout ;
wire \Mux15~13_combout ;
wire \Mux15~16_combout ;
wire \Mux15~19_combout ;
wire \Mux15~7_combout ;
wire \Mux15~8_combout ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \regs[26][16]~q ;
wire \Mux15~2_combout ;
wire \Mux15~3_combout ;
wire \Mux15~6_combout ;
wire \Mux15~9_combout ;
wire \regs~31_combout ;
wire \regs~32_combout ;
wire \regs[26][15]~q ;
wire \regs[30][15]~q ;
wire \regs[22][15]~q ;
wire \regs[18][15]~q ;
wire \Mux48~2_combout ;
wire \Mux48~3_combout ;
wire \regs[20][15]~q ;
wire \regs[16][15]~feeder_combout ;
wire \regs[16][15]~q ;
wire \Mux48~4_combout ;
wire \regs[28][15]~q ;
wire \Mux48~5_combout ;
wire \Mux48~6_combout ;
wire \regs[21][15]~q ;
wire \regs[29][15]~q ;
wire \regs[25][15]~feeder_combout ;
wire \regs[25][15]~q ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \regs[23][15]~q ;
wire \regs[31][15]~q ;
wire \regs[27][15]~feeder_combout ;
wire \regs[27][15]~q ;
wire \regs[19][15]~q ;
wire \Mux48~7_combout ;
wire \Mux48~8_combout ;
wire \regs[6][15]~q ;
wire \regs[7][15]~q ;
wire \regs[4][15]~q ;
wire \regs[5][15]~q ;
wire \Mux48~10_combout ;
wire \Mux48~11_combout ;
wire \regs[15][15]~feeder_combout ;
wire \regs[15][15]~q ;
wire \regs[14][15]~q ;
wire \regs[12][15]~q ;
wire \Mux48~17_combout ;
wire \Mux48~18_combout ;
wire \regs[2][15]~q ;
wire \regs[1][15]~q ;
wire \Mux48~14_combout ;
wire \Mux48~15_combout ;
wire \regs[9][15]~feeder_combout ;
wire \regs[9][15]~q ;
wire \regs[11][15]~q ;
wire \regs[8][15]~q ;
wire \Mux48~12_combout ;
wire \Mux48~13_combout ;
wire \Mux48~16_combout ;
wire \regs[3][15]~q ;
wire \Mux16~14_combout ;
wire \Mux16~15_combout ;
wire \Mux16~12_combout ;
wire \Mux16~13_combout ;
wire \Mux16~16_combout ;
wire \Mux16~18_combout ;
wire \regs[10][15]~q ;
wire \Mux16~10_combout ;
wire \Mux16~11_combout ;
wire \Mux16~19_combout ;
wire \Mux16~8_combout ;
wire \regs[24][15]~q ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~6_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux16~9_combout ;
wire \regs~33_combout ;
wire \regs~34_combout ;
wire \regs[29][14]~feeder_combout ;
wire \regs[29][14]~q ;
wire \regs[25][14]~q ;
wire \regs[21][14]~feeder_combout ;
wire \regs[21][14]~q ;
wire \regs[17][14]~q ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \regs[20][14]~q ;
wire \regs[28][14]~q ;
wire \regs[24][14]~feeder_combout ;
wire \regs[24][14]~q ;
wire \regs[16][14]~q ;
wire \Mux49~4_combout ;
wire \Mux49~5_combout ;
wire \regs[30][14]~q ;
wire \regs[18][14]~q ;
wire \Mux49~2_combout ;
wire \Mux49~3_combout ;
wire \Mux49~6_combout ;
wire \regs[27][14]~q ;
wire \regs[31][14]~q ;
wire \regs[23][14]~q ;
wire \regs[19][14]~q ;
wire \Mux49~7_combout ;
wire \Mux49~8_combout ;
wire \regs[9][14]~q ;
wire \regs[11][14]~q ;
wire \regs[10][14]~q ;
wire \regs[8][14]~q ;
wire \Mux49~10_combout ;
wire \Mux49~11_combout ;
wire \regs[15][14]~feeder_combout ;
wire \regs[15][14]~q ;
wire \regs[14][14]~q ;
wire \regs[12][14]~feeder_combout ;
wire \regs[12][14]~q ;
wire \Mux49~17_combout ;
wire \Mux49~18_combout ;
wire \regs[6][14]~q ;
wire \regs[7][14]~q ;
wire \Mux49~13_combout ;
wire \regs[2][14]~q ;
wire \regs[1][14]~q ;
wire \regs[3][14]~q ;
wire \Mux49~14_combout ;
wire \Mux49~15_combout ;
wire \Mux49~16_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Mux17~7_combout ;
wire \Mux17~8_combout ;
wire \Mux17~4_combout ;
wire \Mux17~5_combout ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux17~6_combout ;
wire \Mux17~9_combout ;
wire \Mux17~14_combout ;
wire \Mux17~15_combout ;
wire \Mux17~12_combout ;
wire \Mux17~13_combout ;
wire \Mux17~16_combout ;
wire \Mux17~18_combout ;
wire \regs[4][14]~q ;
wire \regs[5][14]~q ;
wire \Mux17~10_combout ;
wire \Mux17~11_combout ;
wire \Mux17~19_combout ;
wire \regs~35_combout ;
wire \regs~36_combout ;
wire \regs[23][13]~q ;
wire \regs[31][13]~q ;
wire \regs[19][13]~feeder_combout ;
wire \regs[19][13]~q ;
wire \Mux50~7_combout ;
wire \Mux50~8_combout ;
wire \regs[18][13]~q ;
wire \Mux50~2_combout ;
wire \regs[30][13]~q ;
wire \Mux50~3_combout ;
wire \regs[24][13]~q ;
wire \regs[28][13]~q ;
wire \regs[16][13]~q ;
wire \Mux50~4_combout ;
wire \Mux50~5_combout ;
wire \Mux50~6_combout ;
wire \regs[21][13]~q ;
wire \regs[29][13]~feeder_combout ;
wire \regs[29][13]~q ;
wire \regs[25][13]~q ;
wire \regs[17][13]~q ;
wire \Mux50~0_combout ;
wire \Mux50~1_combout ;
wire \regs[15][13]~feeder_combout ;
wire \regs[15][13]~q ;
wire \regs[14][13]~q ;
wire \regs[13][13]~q ;
wire \Mux50~17_combout ;
wire \Mux50~18_combout ;
wire \regs[6][13]~q ;
wire \regs[7][13]~q ;
wire \regs[5][13]~q ;
wire \regs[4][13]~q ;
wire \Mux50~10_combout ;
wire \Mux50~11_combout ;
wire \regs[9][13]~feeder_combout ;
wire \regs[9][13]~q ;
wire \regs[11][13]~q ;
wire \regs[10][13]~q ;
wire \regs[8][13]~q ;
wire \Mux50~12_combout ;
wire \Mux50~13_combout ;
wire \regs[2][13]~q ;
wire \regs[1][13]~q ;
wire \Mux50~14_combout ;
wire \Mux50~15_combout ;
wire \Mux50~16_combout ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \regs[20][13]~q ;
wire \Mux18~4_combout ;
wire \Mux18~5_combout ;
wire \regs[22][13]~q ;
wire \regs[26][13]~q ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \Mux18~6_combout ;
wire \regs[27][13]~q ;
wire \Mux18~7_combout ;
wire \Mux18~8_combout ;
wire \Mux18~9_combout ;
wire \regs[12][13]~feeder_combout ;
wire \regs[12][13]~q ;
wire \Mux18~17_combout ;
wire \Mux18~18_combout ;
wire \Mux18~10_combout ;
wire \Mux18~11_combout ;
wire \Mux18~12_combout ;
wire \Mux18~13_combout ;
wire \Mux18~14_combout ;
wire \Mux18~15_combout ;
wire \Mux18~16_combout ;
wire \Mux18~19_combout ;
wire \regs~37_combout ;
wire \regs~38_combout ;
wire \regs[31][12]~feeder_combout ;
wire \regs[31][12]~q ;
wire \regs[27][12]~q ;
wire \regs[19][12]~q ;
wire \regs[23][12]~q ;
wire \Mux51~7_combout ;
wire \Mux51~8_combout ;
wire \regs[21][12]~q ;
wire \regs[17][12]~q ;
wire \Mux51~0_combout ;
wire \regs[25][12]~q ;
wire \regs[29][12]~q ;
wire \Mux51~1_combout ;
wire \regs[20][12]~q ;
wire \regs[28][12]~q ;
wire \regs[16][12]~q ;
wire \Mux51~4_combout ;
wire \Mux51~5_combout ;
wire \regs[30][12]~q ;
wire \regs[18][12]~q ;
wire \Mux51~2_combout ;
wire \Mux51~3_combout ;
wire \Mux51~6_combout ;
wire \regs[8][12]~q ;
wire \regs[10][12]~q ;
wire \Mux51~10_combout ;
wire \regs[11][12]~q ;
wire \regs[9][12]~q ;
wire \Mux51~11_combout ;
wire \regs[14][12]~feeder_combout ;
wire \regs[14][12]~q ;
wire \regs[15][12]~q ;
wire \regs[13][12]~q ;
wire \regs[12][12]~q ;
wire \Mux51~17_combout ;
wire \Mux51~18_combout ;
wire \regs[6][12]~q ;
wire \regs[7][12]~q ;
wire \regs[4][12]~q ;
wire \Mux51~12_combout ;
wire \Mux51~13_combout ;
wire \regs[2][12]~q ;
wire \regs[1][12]~q ;
wire \Mux51~14_combout ;
wire \Mux51~15_combout ;
wire \Mux51~16_combout ;
wire \Mux19~1_combout ;
wire \regs[26][12]~feeder_combout ;
wire \regs[26][12]~q ;
wire \regs[22][12]~q ;
wire \Mux19~2_combout ;
wire \Mux19~3_combout ;
wire \Mux19~4_combout ;
wire \Mux19~5_combout ;
wire \Mux19~6_combout ;
wire \Mux19~7_combout ;
wire \Mux19~8_combout ;
wire \Mux19~9_combout ;
wire \regs[5][12]~q ;
wire \Mux19~10_combout ;
wire \Mux19~11_combout ;
wire \Mux19~17_combout ;
wire \Mux19~18_combout ;
wire \Mux19~12_combout ;
wire \Mux19~13_combout ;
wire \regs[3][12]~q ;
wire \Mux19~14_combout ;
wire \Mux19~15_combout ;
wire \Mux19~16_combout ;
wire \Mux19~19_combout ;
wire \regs~39_combout ;
wire \regs~40_combout ;
wire \regs[23][11]~feeder_combout ;
wire \regs[23][11]~q ;
wire \regs[19][11]~q ;
wire \regs[27][11]~q ;
wire \Mux52~7_combout ;
wire \regs[31][11]~q ;
wire \Mux52~8_combout ;
wire \regs[29][11]~q ;
wire \regs[21][11]~feeder_combout ;
wire \regs[21][11]~q ;
wire \regs[25][11]~feeder_combout ;
wire \regs[25][11]~q ;
wire \Mux52~0_combout ;
wire \Mux52~1_combout ;
wire \regs[20][11]~q ;
wire \Mux52~4_combout ;
wire \regs[24][11]~q ;
wire \Mux52~5_combout ;
wire \regs[26][11]~feeder_combout ;
wire \regs[26][11]~q ;
wire \regs[22][11]~q ;
wire \Mux52~2_combout ;
wire \Mux52~3_combout ;
wire \Mux52~6_combout ;
wire \regs[14][11]~q ;
wire \regs[15][11]~feeder_combout ;
wire \regs[15][11]~q ;
wire \regs[12][11]~q ;
wire \Mux52~17_combout ;
wire \Mux52~18_combout ;
wire \regs[2][11]~q ;
wire \regs[3][11]~q ;
wire \regs[1][11]~q ;
wire \Mux52~14_combout ;
wire \Mux52~15_combout ;
wire \regs[9][11]~feeder_combout ;
wire \regs[9][11]~q ;
wire \regs[11][11]~q ;
wire \regs[10][11]~q ;
wire \regs[8][11]~q ;
wire \Mux52~12_combout ;
wire \Mux52~13_combout ;
wire \Mux52~16_combout ;
wire \regs[7][11]~q ;
wire \regs[5][11]~q ;
wire \Mux52~10_combout ;
wire \regs[6][11]~q ;
wire \Mux52~11_combout ;
wire \regs[4][11]~q ;
wire \Mux20~12_combout ;
wire \Mux20~13_combout ;
wire \Mux20~14_combout ;
wire \Mux20~15_combout ;
wire \Mux20~16_combout ;
wire \Mux20~18_combout ;
wire \Mux20~10_combout ;
wire \Mux20~11_combout ;
wire \Mux20~19_combout ;
wire \Mux20~7_combout ;
wire \Mux20~8_combout ;
wire \regs[17][11]~feeder_combout ;
wire \regs[17][11]~q ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \regs[28][11]~q ;
wire \regs[16][11]~q ;
wire \Mux20~4_combout ;
wire \Mux20~5_combout ;
wire \regs[18][11]~feeder_combout ;
wire \regs[18][11]~q ;
wire \Mux20~2_combout ;
wire \Mux20~3_combout ;
wire \Mux20~6_combout ;
wire \Mux20~9_combout ;
wire \regs~41_combout ;
wire \regs~42_combout ;
wire \regs[27][10]~q ;
wire \regs[31][10]~q ;
wire \regs[19][10]~feeder_combout ;
wire \regs[19][10]~q ;
wire \Mux53~7_combout ;
wire \Mux53~8_combout ;
wire \regs[30][10]~q ;
wire \regs[18][10]~q ;
wire \Mux53~2_combout ;
wire \Mux53~3_combout ;
wire \regs[28][10]~q ;
wire \regs[20][10]~q ;
wire \regs[24][10]~q ;
wire \Mux53~4_combout ;
wire \Mux53~5_combout ;
wire \Mux53~6_combout ;
wire \regs[29][10]~feeder_combout ;
wire \regs[29][10]~q ;
wire \regs[25][10]~q ;
wire \regs[21][10]~q ;
wire \Mux53~0_combout ;
wire \Mux53~1_combout ;
wire \regs[14][10]~q ;
wire \regs[15][10]~q ;
wire \regs[13][10]~q ;
wire \regs[12][10]~q ;
wire \Mux53~17_combout ;
wire \Mux53~18_combout ;
wire \regs[11][10]~q ;
wire \regs[10][10]~q ;
wire \Mux53~10_combout ;
wire \regs[9][10]~q ;
wire \Mux53~11_combout ;
wire \regs[2][10]~q ;
wire \regs[1][10]~q ;
wire \Mux53~14_combout ;
wire \Mux53~15_combout ;
wire \regs[7][10]~q ;
wire \regs[5][10]~feeder_combout ;
wire \regs[5][10]~q ;
wire \regs[4][10]~q ;
wire \Mux53~12_combout ;
wire \Mux53~13_combout ;
wire \Mux53~16_combout ;
wire \regs[23][10]~q ;
wire \Mux21~7_combout ;
wire \Mux21~8_combout ;
wire \regs[16][10]~feeder_combout ;
wire \regs[16][10]~q ;
wire \Mux21~4_combout ;
wire \Mux21~5_combout ;
wire \Mux21~6_combout ;
wire \regs[17][10]~q ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux21~9_combout ;
wire \regs[6][10]~feeder_combout ;
wire \regs[6][10]~q ;
wire \Mux21~10_combout ;
wire \Mux21~11_combout ;
wire \Mux21~17_combout ;
wire \Mux21~18_combout ;
wire \regs[8][10]~q ;
wire \Mux21~12_combout ;
wire \Mux21~13_combout ;
wire \regs[3][10]~feeder_combout ;
wire \regs[3][10]~q ;
wire \Mux21~14_combout ;
wire \Mux21~15_combout ;
wire \Mux21~16_combout ;
wire \Mux21~19_combout ;
wire \regs~43_combout ;
wire \regs~44_combout ;
wire \regs[29][9]~feeder_combout ;
wire \regs[29][9]~q ;
wire \regs[21][9]~feeder_combout ;
wire \regs[21][9]~q ;
wire \regs[17][9]~q ;
wire \regs[25][9]~q ;
wire \Mux54~0_combout ;
wire \Mux54~1_combout ;
wire \regs[24][9]~q ;
wire \regs[20][9]~q ;
wire \Mux54~4_combout ;
wire \Mux54~5_combout ;
wire \regs[30][9]~feeder_combout ;
wire \regs[30][9]~q ;
wire \regs[26][9]~q ;
wire \regs[18][9]~q ;
wire \regs[22][9]~q ;
wire \Mux54~2_combout ;
wire \Mux54~3_combout ;
wire \Mux54~6_combout ;
wire \regs[31][9]~q ;
wire \regs[23][9]~q ;
wire \regs[27][9]~feeder_combout ;
wire \regs[27][9]~q ;
wire \Mux54~7_combout ;
wire \Mux54~8_combout ;
wire \regs[15][9]~q ;
wire \regs[14][9]~feeder_combout ;
wire \regs[14][9]~q ;
wire \regs[13][9]~q ;
wire \regs[12][9]~q ;
wire \Mux54~17_combout ;
wire \Mux54~18_combout ;
wire \regs[5][9]~q ;
wire \Mux54~10_combout ;
wire \regs[7][9]~q ;
wire \regs[6][9]~q ;
wire \Mux54~11_combout ;
wire \regs[9][9]~q ;
wire \regs[11][9]~q ;
wire \regs[10][9]~q ;
wire \regs[8][9]~q ;
wire \Mux54~12_combout ;
wire \Mux54~13_combout ;
wire \regs[2][9]~q ;
wire \regs[1][9]~q ;
wire \Mux54~14_combout ;
wire \Mux54~15_combout ;
wire \Mux54~16_combout ;
wire \regs[19][9]~q ;
wire \Mux22~7_combout ;
wire \Mux22~8_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \regs[16][9]~feeder_combout ;
wire \regs[16][9]~q ;
wire \Mux22~4_combout ;
wire \Mux22~5_combout ;
wire \Mux22~2_combout ;
wire \Mux22~3_combout ;
wire \Mux22~6_combout ;
wire \Mux22~9_combout ;
wire \Mux22~11_combout ;
wire \Mux22~17_combout ;
wire \Mux22~18_combout ;
wire \regs[3][9]~feeder_combout ;
wire \regs[3][9]~q ;
wire \Mux22~14_combout ;
wire \Mux22~15_combout ;
wire \regs[4][9]~q ;
wire \Mux22~12_combout ;
wire \Mux22~13_combout ;
wire \Mux22~16_combout ;
wire \Mux22~19_combout ;
wire \regs~45_combout ;
wire \regs~46_combout ;
wire \regs[22][8]~q ;
wire \regs[30][8]~q ;
wire \Mux55~3_combout ;
wire \regs[20][8]~q ;
wire \regs[24][8]~q ;
wire \Mux55~4_combout ;
wire \Mux55~5_combout ;
wire \Mux55~6_combout ;
wire \regs[29][8]~feeder_combout ;
wire \regs[29][8]~q ;
wire \regs[25][8]~q ;
wire \regs[17][8]~q ;
wire \Mux55~0_combout ;
wire \Mux55~1_combout ;
wire \regs[31][8]~q ;
wire \regs[27][8]~q ;
wire \regs[19][8]~q ;
wire \Mux55~7_combout ;
wire \Mux55~8_combout ;
wire \regs[11][8]~q ;
wire \regs[9][8]~q ;
wire \regs[10][8]~q ;
wire \Mux55~10_combout ;
wire \Mux55~11_combout ;
wire \regs[15][8]~q ;
wire \regs[14][8]~q ;
wire \regs[12][8]~q ;
wire \Mux55~17_combout ;
wire \Mux55~18_combout ;
wire \regs[2][8]~q ;
wire \regs[3][8]~feeder_combout ;
wire \regs[3][8]~q ;
wire \regs[1][8]~q ;
wire \Mux55~14_combout ;
wire \Mux55~15_combout ;
wire \regs[6][8]~q ;
wire \regs[7][8]~q ;
wire \regs[5][8]~q ;
wire \regs[4][8]~q ;
wire \Mux55~12_combout ;
wire \Mux55~13_combout ;
wire \Mux55~16_combout ;
wire \regs[18][8]~q ;
wire \Mux23~2_combout ;
wire \Mux23~3_combout ;
wire \regs[28][8]~q ;
wire \regs[16][8]~q ;
wire \Mux23~4_combout ;
wire \Mux23~5_combout ;
wire \Mux23~6_combout ;
wire \regs[21][8]~feeder_combout ;
wire \regs[21][8]~q ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \Mux23~7_combout ;
wire \Mux23~8_combout ;
wire \Mux23~9_combout ;
wire \regs[13][8]~feeder_combout ;
wire \regs[13][8]~q ;
wire \Mux23~17_combout ;
wire \Mux23~18_combout ;
wire \Mux23~10_combout ;
wire \Mux23~11_combout ;
wire \regs[8][8]~q ;
wire \Mux23~12_combout ;
wire \Mux23~13_combout ;
wire \Mux23~14_combout ;
wire \Mux23~15_combout ;
wire \Mux23~16_combout ;
wire \Mux23~19_combout ;
wire \regs~47_combout ;
wire \regs~48_combout ;
wire \regs~49_combout ;
wire \regs[21][7]~q ;
wire \regs[29][7]~q ;
wire \regs[17][7]~q ;
wire \regs[25][7]~q ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \regs[30][7]~feeder_combout ;
wire \regs[30][7]~q ;
wire \regs[26][7]~q ;
wire \Mux56~3_combout ;
wire \regs[24][7]~q ;
wire \regs[20][7]~q ;
wire \Mux56~4_combout ;
wire \Mux56~5_combout ;
wire \Mux56~6_combout ;
wire \regs[31][7]~q ;
wire \regs[23][7]~q ;
wire \regs[19][7]~feeder_combout ;
wire \regs[19][7]~q ;
wire \regs[27][7]~q ;
wire \Mux56~7_combout ;
wire \Mux56~8_combout ;
wire \regs[14][7]~q ;
wire \regs[15][7]~q ;
wire \regs[13][7]~feeder_combout ;
wire \regs[13][7]~q ;
wire \regs[12][7]~q ;
wire \Mux56~17_combout ;
wire \Mux56~18_combout ;
wire \regs[7][7]~q ;
wire \regs[6][7]~q ;
wire \regs[5][7]~q ;
wire \Mux56~10_combout ;
wire \Mux56~11_combout ;
wire \regs[10][7]~q ;
wire \regs[8][7]~q ;
wire \Mux56~12_combout ;
wire \regs[11][7]~q ;
wire \regs[9][7]~q ;
wire \Mux56~13_combout ;
wire \regs[2][7]~q ;
wire \regs[1][7]~q ;
wire \Mux56~14_combout ;
wire \Mux56~15_combout ;
wire \Mux56~16_combout ;
wire \Mux24~10_combout ;
wire \Mux24~11_combout ;
wire \Mux24~17_combout ;
wire \Mux24~18_combout ;
wire \regs[4][7]~q ;
wire \Mux24~12_combout ;
wire \Mux24~13_combout ;
wire \regs[3][7]~q ;
wire \Mux24~14_combout ;
wire \Mux24~15_combout ;
wire \Mux24~16_combout ;
wire \Mux24~19_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \regs[28][7]~q ;
wire \regs[16][7]~q ;
wire \Mux24~4_combout ;
wire \Mux24~5_combout ;
wire \regs[22][7]~q ;
wire \regs[18][7]~feeder_combout ;
wire \regs[18][7]~q ;
wire \Mux24~2_combout ;
wire \Mux24~3_combout ;
wire \Mux24~6_combout ;
wire \Mux24~7_combout ;
wire \Mux24~8_combout ;
wire \Mux24~9_combout ;
wire \regs~50_combout ;
wire \regs~51_combout ;
wire \regs~52_combout ;
wire \regs[25][6]~q ;
wire \regs[29][6]~feeder_combout ;
wire \regs[29][6]~q ;
wire \regs[21][6]~q ;
wire \Mux57~0_combout ;
wire \Mux57~1_combout ;
wire \regs[31][6]~q ;
wire \regs[27][6]~feeder_combout ;
wire \regs[27][6]~q ;
wire \regs[23][6]~feeder_combout ;
wire \regs[23][6]~q ;
wire \Mux57~7_combout ;
wire \Mux57~8_combout ;
wire \regs[22][6]~q ;
wire \regs[30][6]~q ;
wire \Mux57~3_combout ;
wire \regs[28][6]~q ;
wire \regs[20][6]~q ;
wire \regs[16][6]~q ;
wire \regs[24][6]~q ;
wire \Mux57~4_combout ;
wire \Mux57~5_combout ;
wire \Mux57~6_combout ;
wire \regs[14][6]~q ;
wire \regs[15][6]~q ;
wire \regs[13][6]~q ;
wire \regs[12][6]~q ;
wire \Mux57~17_combout ;
wire \Mux57~18_combout ;
wire \regs[11][6]~q ;
wire \regs[9][6]~q ;
wire \regs[10][6]~q ;
wire \Mux57~10_combout ;
wire \Mux57~11_combout ;
wire \regs[2][6]~q ;
wire \regs[3][6]~q ;
wire \regs[1][6]~q ;
wire \Mux57~14_combout ;
wire \Mux57~15_combout ;
wire \regs[6][6]~feeder_combout ;
wire \regs[6][6]~q ;
wire \regs[7][6]~q ;
wire \regs[4][6]~q ;
wire \Mux57~12_combout ;
wire \Mux57~13_combout ;
wire \Mux57~16_combout ;
wire \regs[19][6]~q ;
wire \Mux25~7_combout ;
wire \Mux25~8_combout ;
wire \regs[18][6]~q ;
wire \Mux25~2_combout ;
wire \Mux25~3_combout ;
wire \Mux25~4_combout ;
wire \Mux25~5_combout ;
wire \Mux25~6_combout ;
wire \regs[17][6]~feeder_combout ;
wire \regs[17][6]~q ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux25~9_combout ;
wire \regs[5][6]~q ;
wire \Mux25~10_combout ;
wire \Mux25~11_combout ;
wire \Mux25~17_combout ;
wire \Mux25~18_combout ;
wire \Mux25~14_combout ;
wire \Mux25~15_combout ;
wire \Mux25~12_combout ;
wire \Mux25~13_combout ;
wire \Mux25~16_combout ;
wire \Mux25~19_combout ;
wire \regs~53_combout ;
wire \regs~54_combout ;
wire \regs~55_combout ;
wire \regs[23][5]~feeder_combout ;
wire \regs[23][5]~q ;
wire \regs[27][5]~feeder_combout ;
wire \regs[27][5]~q ;
wire \Mux58~7_combout ;
wire \regs[31][5]~q ;
wire \Mux58~8_combout ;
wire \regs[21][5]~feeder_combout ;
wire \regs[21][5]~q ;
wire \regs[29][5]~feeder_combout ;
wire \regs[29][5]~q ;
wire \regs[25][5]~feeder_combout ;
wire \regs[25][5]~q ;
wire \Mux58~0_combout ;
wire \Mux58~1_combout ;
wire \regs[22][5]~q ;
wire \Mux58~2_combout ;
wire \regs[26][5]~q ;
wire \Mux58~3_combout ;
wire \regs[24][5]~feeder_combout ;
wire \regs[24][5]~q ;
wire \regs[20][5]~feeder_combout ;
wire \regs[20][5]~q ;
wire \Mux58~4_combout ;
wire \Mux58~5_combout ;
wire \Mux58~6_combout ;
wire \regs[14][5]~q ;
wire \regs[15][5]~q ;
wire \regs[12][5]~q ;
wire \Mux58~17_combout ;
wire \Mux58~18_combout ;
wire \regs[9][5]~feeder_combout ;
wire \regs[9][5]~q ;
wire \regs[11][5]~q ;
wire \regs[10][5]~q ;
wire \regs[8][5]~q ;
wire \Mux58~12_combout ;
wire \Mux58~13_combout ;
wire \regs[2][5]~feeder_combout ;
wire \regs[2][5]~q ;
wire \regs[1][5]~q ;
wire \Mux58~14_combout ;
wire \Mux58~15_combout ;
wire \Mux58~16_combout ;
wire \regs[7][5]~q ;
wire \regs[6][5]~q ;
wire \regs[5][5]~q ;
wire \Mux58~10_combout ;
wire \Mux58~11_combout ;
wire \Mux26~10_combout ;
wire \Mux26~11_combout ;
wire \regs[3][5]~q ;
wire \Mux26~14_combout ;
wire \Mux26~15_combout ;
wire \regs[4][5]~q ;
wire \Mux26~12_combout ;
wire \Mux26~13_combout ;
wire \Mux26~16_combout ;
wire \regs[13][5]~q ;
wire \Mux26~17_combout ;
wire \Mux26~18_combout ;
wire \Mux26~19_combout ;
wire \Mux26~1_combout ;
wire \Mux26~8_combout ;
wire \regs[28][5]~q ;
wire \regs[16][5]~feeder_combout ;
wire \regs[16][5]~q ;
wire \Mux26~4_combout ;
wire \Mux26~5_combout ;
wire \Mux26~2_combout ;
wire \Mux26~3_combout ;
wire \Mux26~6_combout ;
wire \Mux26~9_combout ;
wire \regs~56_combout ;
wire \regs~57_combout ;
wire \regs~58_combout ;
wire \regs[27][4]~feeder_combout ;
wire \regs[27][4]~q ;
wire \regs[31][4]~q ;
wire \regs[23][4]~feeder_combout ;
wire \regs[23][4]~q ;
wire \regs[19][4]~q ;
wire \Mux59~7_combout ;
wire \Mux59~8_combout ;
wire \regs[22][4]~q ;
wire \regs[26][4]~q ;
wire \Mux59~2_combout ;
wire \Mux59~3_combout ;
wire \regs[28][4]~q ;
wire \regs[20][4]~q ;
wire \Mux59~5_combout ;
wire \Mux59~6_combout ;
wire \regs[25][4]~q ;
wire \regs[29][4]~q ;
wire \regs[21][4]~q ;
wire \Mux59~0_combout ;
wire \Mux59~1_combout ;
wire \regs[15][4]~q ;
wire \regs[14][4]~q ;
wire \regs[12][4]~q ;
wire \regs[13][4]~q ;
wire \Mux59~17_combout ;
wire \Mux59~18_combout ;
wire \regs[10][4]~q ;
wire \Mux59~10_combout ;
wire \regs[11][4]~q ;
wire \regs[9][4]~q ;
wire \Mux59~11_combout ;
wire \regs[1][4]~q ;
wire \regs[3][4]~q ;
wire \Mux59~14_combout ;
wire \regs[2][4]~q ;
wire \Mux59~15_combout ;
wire \regs[7][4]~q ;
wire \regs[6][4]~q ;
wire \Mux59~13_combout ;
wire \Mux59~16_combout ;
wire \regs[30][4]~q ;
wire \regs[18][4]~q ;
wire \Mux27~2_combout ;
wire \Mux27~3_combout ;
wire \Mux27~6_combout ;
wire \Mux27~7_combout ;
wire \Mux27~8_combout ;
wire \regs[17][4]~q ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Mux27~9_combout ;
wire \Mux27~17_combout ;
wire \Mux27~18_combout ;
wire \regs[4][4]~q ;
wire \regs[5][4]~q ;
wire \Mux27~10_combout ;
wire \Mux27~11_combout ;
wire \regs[8][4]~q ;
wire \Mux27~12_combout ;
wire \Mux27~13_combout ;
wire \Mux27~16_combout ;
wire \Mux27~19_combout ;
wire \regs~60_combout ;
wire \regs[29][3]~q ;
wire \regs[17][3]~feeder_combout ;
wire \regs[17][3]~q ;
wire \regs[25][3]~q ;
wire \Mux60~0_combout ;
wire \regs[21][3]~q ;
wire \Mux60~1_combout ;
wire \regs[30][3]~q ;
wire \regs[26][3]~q ;
wire \regs[22][3]~q ;
wire \Mux60~2_combout ;
wire \Mux60~3_combout ;
wire \regs[28][3]~q ;
wire \regs[24][3]~q ;
wire \Mux60~5_combout ;
wire \Mux60~6_combout ;
wire \regs[23][3]~feeder_combout ;
wire \regs[23][3]~q ;
wire \regs[31][3]~q ;
wire \regs[19][3]~q ;
wire \Mux60~7_combout ;
wire \Mux60~8_combout ;
wire \regs[14][3]~feeder_combout ;
wire \regs[14][3]~q ;
wire \regs[13][3]~q ;
wire \Mux60~17_combout ;
wire \regs[15][3]~q ;
wire \Mux60~18_combout ;
wire \regs[7][3]~q ;
wire \regs[6][3]~q ;
wire \regs[5][3]~q ;
wire \Mux60~10_combout ;
wire \Mux60~11_combout ;
wire \regs[2][3]~q ;
wire \regs[3][3]~q ;
wire \regs[1][3]~q ;
wire \Mux60~14_combout ;
wire \Mux60~15_combout ;
wire \regs[11][3]~q ;
wire \regs[9][3]~q ;
wire \regs[8][3]~feeder_combout ;
wire \regs[8][3]~q ;
wire \Mux60~12_combout ;
wire \Mux60~13_combout ;
wire \Mux60~16_combout ;
wire \Mux28~7_combout ;
wire \Mux28~8_combout ;
wire \regs[18][3]~feeder_combout ;
wire \regs[18][3]~q ;
wire \Mux28~2_combout ;
wire \Mux28~3_combout ;
wire \regs[20][3]~q ;
wire \regs[16][3]~q ;
wire \Mux28~4_combout ;
wire \Mux28~5_combout ;
wire \Mux28~6_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Mux28~9_combout ;
wire \regs[10][3]~feeder_combout ;
wire \regs[10][3]~q ;
wire \Mux28~10_combout ;
wire \Mux28~11_combout ;
wire \regs[12][3]~q ;
wire \Mux28~17_combout ;
wire \Mux28~18_combout ;
wire \regs[4][3]~q ;
wire \Mux28~12_combout ;
wire \Mux28~13_combout ;
wire \Mux28~16_combout ;
wire \Mux28~19_combout ;
wire \regs~61_combout ;
wire \regs~62_combout ;
wire \regs[20][2]~q ;
wire \regs[16][2]~q ;
wire \regs[24][2]~q ;
wire \Mux61~4_combout ;
wire \Mux61~5_combout ;
wire \regs[22][2]~q ;
wire \regs[26][2]~q ;
wire \Mux61~2_combout ;
wire \Mux61~3_combout ;
wire \Mux61~6_combout ;
wire \regs[27][2]~feeder_combout ;
wire \regs[27][2]~q ;
wire \regs[23][2]~feeder_combout ;
wire \regs[23][2]~q ;
wire \regs[19][2]~q ;
wire \Mux61~7_combout ;
wire \regs[31][2]~q ;
wire \Mux61~8_combout ;
wire \regs[29][2]~q ;
wire \regs[25][2]~feeder_combout ;
wire \regs[25][2]~q ;
wire \regs[17][2]~feeder_combout ;
wire \regs[17][2]~q ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \regs[15][2]~q ;
wire \regs[14][2]~q ;
wire \regs[13][2]~q ;
wire \Mux61~17_combout ;
wire \Mux61~18_combout ;
wire \regs[2][2]~q ;
wire \regs[3][2]~feeder_combout ;
wire \regs[3][2]~q ;
wire \Mux61~14_combout ;
wire \Mux61~15_combout ;
wire \regs[6][2]~q ;
wire \regs[7][2]~q ;
wire \regs[4][2]~q ;
wire \Mux61~12_combout ;
wire \Mux61~13_combout ;
wire \Mux61~16_combout ;
wire \regs[9][2]~feeder_combout ;
wire \regs[9][2]~q ;
wire \regs[11][2]~feeder_combout ;
wire \regs[11][2]~q ;
wire \regs[10][2]~feeder_combout ;
wire \regs[10][2]~q ;
wire \Mux61~10_combout ;
wire \Mux61~11_combout ;
wire \regs[28][2]~q ;
wire \Mux29~4_combout ;
wire \Mux29~5_combout ;
wire \regs[30][2]~q ;
wire \regs[18][2]~q ;
wire \Mux29~2_combout ;
wire \Mux29~3_combout ;
wire \Mux29~6_combout ;
wire \Mux29~7_combout ;
wire \Mux29~8_combout ;
wire \regs[21][2]~feeder_combout ;
wire \regs[21][2]~q ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Mux29~9_combout ;
wire \regs[12][2]~q ;
wire \Mux29~17_combout ;
wire \Mux29~18_combout ;
wire \regs[5][2]~q ;
wire \Mux29~10_combout ;
wire \Mux29~11_combout ;
wire \regs[1][2]~q ;
wire \Mux29~14_combout ;
wire \Mux29~15_combout ;
wire \regs[8][2]~q ;
wire \Mux29~12_combout ;
wire \Mux29~13_combout ;
wire \Mux29~16_combout ;
wire \Mux29~19_combout ;
wire \regs[16][1]~q ;
wire \Mux62~4_combout ;
wire \Mux62~5_combout ;
wire \regs[30][1]~q ;
wire \Mux62~2_combout ;
wire \Mux62~3_combout ;
wire \Mux62~6_combout ;
wire \regs[17][1]~q ;
wire \Mux62~0_combout ;
wire \Mux62~1_combout ;
wire \regs[23][1]~feeder_combout ;
wire \regs[23][1]~q ;
wire \Mux62~7_combout ;
wire \Mux62~8_combout ;
wire \regs[4][1]~q ;
wire \Mux62~10_combout ;
wire \Mux62~11_combout ;
wire \Mux62~17_combout ;
wire \Mux62~18_combout ;
wire \regs[11][1]~q ;
wire \regs[8][1]~q ;
wire \Mux62~12_combout ;
wire \Mux62~13_combout ;
wire \regs[2][1]~q ;
wire \Mux62~14_combout ;
wire \Mux62~15_combout ;
wire \Mux62~16_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \regs[26][0]~feeder_combout ;
wire \regs[26][0]~q ;
wire \Mux31~2_combout ;
wire \Mux31~3_combout ;
wire \Mux31~4_combout ;
wire \Mux31~5_combout ;
wire \Mux31~6_combout ;
wire \regs[19][0]~feeder_combout ;
wire \regs[19][0]~q ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \Mux31~9_combout ;
wire \regs[6][0]~q ;
wire \Mux31~10_combout ;
wire \Mux31~11_combout ;
wire \Mux31~12_combout ;
wire \Mux31~13_combout ;
wire \regs[2][0]~q ;
wire \Mux31~14_combout ;
wire \Mux31~15_combout ;
wire \Mux31~16_combout ;
wire \regs[13][0]~feeder_combout ;
wire \regs[13][0]~q ;
wire \Mux31~17_combout ;
wire \Mux31~18_combout ;
wire \Mux31~19_combout ;
wire \regs~63_combout ;
wire \regs[14][31]~q ;
wire \regs[15][31]~q ;
wire \regs[12][31]~q ;
wire \Mux32~7_combout ;
wire \Mux32~8_combout ;
wire \regs[7][31]~q ;
wire \regs[6][31]~feeder_combout ;
wire \regs[6][31]~q ;
wire \regs[5][31]~feeder_combout ;
wire \regs[5][31]~q ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \regs[2][31]~q ;
wire \regs[1][31]~q ;
wire \Mux32~4_combout ;
wire \Mux32~5_combout ;
wire \regs[9][31]~q ;
wire \regs[11][31]~q ;
wire \regs[10][31]~q ;
wire \regs[8][31]~q ;
wire \Mux32~2_combout ;
wire \Mux32~3_combout ;
wire \Mux32~6_combout ;
wire \regs[31][31]~feeder_combout ;
wire \regs[31][31]~q ;
wire \regs[23][31]~q ;
wire \regs[19][31]~feeder_combout ;
wire \regs[19][31]~q ;
wire \Mux32~17_combout ;
wire \Mux32~18_combout ;
wire \regs[29][31]~feeder_combout ;
wire \regs[29][31]~q ;
wire \regs[21][31]~feeder_combout ;
wire \regs[21][31]~q ;
wire \regs[17][31]~feeder_combout ;
wire \regs[17][31]~q ;
wire \Mux32~10_combout ;
wire \Mux32~11_combout ;
wire \regs[28][31]~q ;
wire \regs[24][31]~q ;
wire \regs[20][31]~q ;
wire \regs[16][31]~q ;
wire \Mux32~14_combout ;
wire \Mux32~15_combout ;
wire \regs[26][31]~feeder_combout ;
wire \regs[26][31]~q ;
wire \regs[18][31]~q ;
wire \regs[22][31]~q ;
wire \Mux32~12_combout ;
wire \Mux32~13_combout ;
wire \Mux32~16_combout ;
wire \regs[13][31]~q ;
wire \Mux0~17_combout ;
wire \Mux0~18_combout ;
wire \Mux0~10_combout ;
wire \Mux0~11_combout ;
wire \regs[3][31]~q ;
wire \Mux0~14_combout ;
wire \Mux0~15_combout ;
wire \Mux0~12_combout ;
wire \Mux0~13_combout ;
wire \Mux0~16_combout ;
wire \Mux0~19_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~7_combout ;
wire \Mux0~8_combout ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \regs[30][31]~q ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~6_combout ;
wire \Mux0~9_combout ;


// Location: FF_X58_Y33_N13
dffeas \regs[21][0] (
	.clk(CLK),
	.d(\regs[21][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][0] .is_wysiwyg = "true";
defparam \regs[21][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N21
dffeas \regs[22][0] (
	.clk(CLK),
	.d(\regs~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][0] .is_wysiwyg = "true";
defparam \regs[22][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N27
dffeas \regs[26][1] (
	.clk(CLK),
	.d(\regs[26][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][1] .is_wysiwyg = "true";
defparam \regs[26][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N11
dffeas \regs[27][1] (
	.clk(CLK),
	.d(\regs[27][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][1] .is_wysiwyg = "true";
defparam \regs[27][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N3
dffeas \regs[1][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][1] .is_wysiwyg = "true";
defparam \regs[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N23
dffeas \regs[17][30] (
	.clk(CLK),
	.d(\regs[17][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][30] .is_wysiwyg = "true";
defparam \regs[17][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N25
dffeas \regs[18][30] (
	.clk(CLK),
	.d(\regs[18][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][30] .is_wysiwyg = "true";
defparam \regs[18][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y43_N31
dffeas \regs[26][29] (
	.clk(CLK),
	.d(\regs[26][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][29] .is_wysiwyg = "true";
defparam \regs[26][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N22
cycloneive_lcell_comb \Mux37~2 (
// Equation(s):
// \Mux37~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[26][26]~q )) # (!dcifimemload_19 & ((\regs[18][26]~q )))))

	.dataa(\regs[26][26]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][26]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux37~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~2 .lut_mask = 16'hEE30;
defparam \Mux37~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N27
dffeas \regs[5][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][26] .is_wysiwyg = "true";
defparam \regs[5][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N26
cycloneive_lcell_comb \Mux5~10 (
// Equation(s):
// \Mux5~10_combout  = (dcifimemload_21 & (((\regs[5][26]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][26]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][26]~q ),
	.datac(\regs[5][26]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux5~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~10 .lut_mask = 16'hAAE4;
defparam \Mux5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N9
dffeas \regs[13][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][25] .is_wysiwyg = "true";
defparam \regs[13][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N22
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\regs[13][25]~q ))) # (!dcifimemload_21 & (\regs[12][25]~q ))))

	.dataa(\regs[12][25]~q ),
	.datab(\regs[13][25]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'hFC0A;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N13
dffeas \regs[18][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][24] .is_wysiwyg = "true";
defparam \regs[18][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N11
dffeas \regs[24][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][24] .is_wysiwyg = "true";
defparam \regs[24][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N10
cycloneive_lcell_comb \Mux39~4 (
// Equation(s):
// \Mux39~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[24][24]~q ))) # (!dcifimemload_19 & (\regs[16][24]~q ))))

	.dataa(\regs[16][24]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[24][24]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux39~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~4 .lut_mask = 16'hFC22;
defparam \Mux39~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N23
dffeas \regs[5][24] (
	.clk(CLK),
	.d(\regs[5][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][24] .is_wysiwyg = "true";
defparam \regs[5][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N12
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (dcifimemload_23 & ((\regs[22][24]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[18][24]~q  & !dcifimemload_24))))

	.dataa(\regs[22][24]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[18][24]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hCCB8;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N25
dffeas \regs[16][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][23] .is_wysiwyg = "true";
defparam \regs[16][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y42_N19
dffeas \regs[28][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][23] .is_wysiwyg = "true";
defparam \regs[28][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N24
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[24][23]~q )) # (!dcifimemload_24 & ((\regs[16][23]~q )))))

	.dataa(\regs[24][23]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[16][23]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'hEE30;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N18
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (dcifimemload_23 & ((\Mux8~4_combout  & ((\regs[28][23]~q ))) # (!\Mux8~4_combout  & (\regs[20][23]~q )))) # (!dcifimemload_23 & (((\Mux8~4_combout ))))

	.dataa(\regs[20][23]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[28][23]~q ),
	.datad(\Mux8~4_combout ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hF388;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N1
dffeas \regs[16][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][22] .is_wysiwyg = "true";
defparam \regs[16][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y45_N31
dffeas \regs[5][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][22] .is_wysiwyg = "true";
defparam \regs[5][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N0
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (dcifimemload_23 & ((\regs[20][22]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[16][22]~q  & !dcifimemload_24))))

	.dataa(\regs[20][22]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[16][22]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hCCB8;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N30
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (dcifimemload_24 & ((\Mux9~4_combout  & ((\regs[28][22]~q ))) # (!\Mux9~4_combout  & (\regs[24][22]~q )))) # (!dcifimemload_24 & (((\Mux9~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[24][22]~q ),
	.datac(\regs[28][22]~q ),
	.datad(\Mux9~4_combout ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hF588;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N30
cycloneive_lcell_comb \Mux9~10 (
// Equation(s):
// \Mux9~10_combout  = (dcifimemload_21 & (((\regs[5][22]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][22]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][22]~q ),
	.datac(\regs[5][22]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~10 .lut_mask = 16'hAAE4;
defparam \Mux9~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N5
dffeas \regs[18][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][21] .is_wysiwyg = "true";
defparam \regs[18][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N4
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[26][21]~q )) # (!dcifimemload_24 & ((\regs[18][21]~q )))))

	.dataa(\regs[26][21]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[18][21]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hEE30;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y32_N27
dffeas \regs[8][19] (
	.clk(CLK),
	.d(\regs[8][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][19] .is_wysiwyg = "true";
defparam \regs[8][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N1
dffeas \regs[26][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][18] .is_wysiwyg = "true";
defparam \regs[26][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N12
cycloneive_lcell_comb \Mux45~4 (
// Equation(s):
// \Mux45~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[24][18]~q )) # (!dcifimemload_19 & ((\regs[16][18]~q )))))

	.dataa(\regs[24][18]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[16][18]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux45~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~4 .lut_mask = 16'hEE30;
defparam \Mux45~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y36_N5
dffeas \regs[3][18] (
	.clk(CLK),
	.d(\regs~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][18] .is_wysiwyg = "true";
defparam \regs[3][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N27
dffeas \regs[13][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][18] .is_wysiwyg = "true";
defparam \regs[13][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N18
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[22][18]~q ))) # (!dcifimemload_23 & (\regs[18][18]~q ))))

	.dataa(dcifimemload_24),
	.datab(\regs[18][18]~q ),
	.datac(\regs[22][18]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hFA44;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N0
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (dcifimemload_24 & ((\Mux13~2_combout  & ((\regs[30][18]~q ))) # (!\Mux13~2_combout  & (\regs[26][18]~q )))) # (!dcifimemload_24 & (\Mux13~2_combout ))

	.dataa(dcifimemload_24),
	.datab(\Mux13~2_combout ),
	.datac(\regs[26][18]~q ),
	.datad(\regs[30][18]~q ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hEC64;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N6
cycloneive_lcell_comb \Mux13~10 (
// Equation(s):
// \Mux13~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\regs[5][18]~q ))) # (!dcifimemload_21 & (\regs[4][18]~q ))))

	.dataa(dcifimemload_22),
	.datab(\regs[4][18]~q ),
	.datac(\regs[5][18]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux13~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~10 .lut_mask = 16'hFA44;
defparam \Mux13~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N26
cycloneive_lcell_comb \Mux13~17 (
// Equation(s):
// \Mux13~17_combout  = (dcifimemload_21 & (((\regs[13][18]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][18]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][18]~q ),
	.datac(\regs[13][18]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux13~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~17 .lut_mask = 16'hAAE4;
defparam \Mux13~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y32_N9
dffeas \regs[8][17] (
	.clk(CLK),
	.d(\regs[8][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][17] .is_wysiwyg = "true";
defparam \regs[8][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N13
dffeas \regs[11][17] (
	.clk(CLK),
	.d(\regs[11][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][17] .is_wysiwyg = "true";
defparam \regs[11][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N13
dffeas \regs[17][15] (
	.clk(CLK),
	.d(\regs[17][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][15] .is_wysiwyg = "true";
defparam \regs[17][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N11
dffeas \regs[13][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][15] .is_wysiwyg = "true";
defparam \regs[13][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N16
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\regs[26][15]~q ))) # (!dcifimemload_24 & (\regs[18][15]~q ))))

	.dataa(dcifimemload_23),
	.datab(\regs[18][15]~q ),
	.datac(\regs[26][15]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hFA44;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N16
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (dcifimemload_23 & ((\Mux16~2_combout  & (\regs[30][15]~q )) # (!\Mux16~2_combout  & ((\regs[22][15]~q ))))) # (!dcifimemload_23 & (((\Mux16~2_combout ))))

	.dataa(\regs[30][15]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[22][15]~q ),
	.datad(\Mux16~2_combout ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hBBC0;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N30
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// \Mux16~7_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\regs[23][15]~q )))) # (!dcifimemload_23 & (!dcifimemload_24 & ((\regs[19][15]~q ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\regs[23][15]~q ),
	.datad(\regs[19][15]~q ),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hB9A8;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N10
cycloneive_lcell_comb \Mux16~17 (
// Equation(s):
// \Mux16~17_combout  = (dcifimemload_21 & (((\regs[13][15]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][15]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][15]~q ),
	.datac(\regs[13][15]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux16~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~17 .lut_mask = 16'hAAE4;
defparam \Mux16~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N11
dffeas \regs[22][14] (
	.clk(CLK),
	.d(\regs[22][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][14] .is_wysiwyg = "true";
defparam \regs[22][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N7
dffeas \regs[26][14] (
	.clk(CLK),
	.d(\regs[26][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][14] .is_wysiwyg = "true";
defparam \regs[26][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N6
cycloneive_lcell_comb \Mux49~12 (
// Equation(s):
// \Mux49~12_combout  = (dcifimemload_16 & ((\regs[5][14]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][14]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[5][14]~q ),
	.datac(\regs[4][14]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux49~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~12 .lut_mask = 16'hAAD8;
defparam \Mux49~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N23
dffeas \regs[13][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][14] .is_wysiwyg = "true";
defparam \regs[13][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N22
cycloneive_lcell_comb \Mux17~17 (
// Equation(s):
// \Mux17~17_combout  = (dcifimemload_21 & (((\regs[13][14]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][14]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][14]~q ),
	.datac(\regs[13][14]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~17 .lut_mask = 16'hAAE4;
defparam \Mux17~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N23
dffeas \regs[3][13] (
	.clk(CLK),
	.d(\regs[3][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][13] .is_wysiwyg = "true";
defparam \regs[3][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N7
dffeas \regs[24][12] (
	.clk(CLK),
	.d(\regs[24][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][12] .is_wysiwyg = "true";
defparam \regs[24][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N10
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (dcifimemload_24 & (((\regs[25][12]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[17][12]~q  & ((!dcifimemload_23))))

	.dataa(\regs[17][12]~q ),
	.datab(\regs[25][12]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hF0CA;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N31
dffeas \regs[30][11] (
	.clk(CLK),
	.d(\regs[30][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][11] .is_wysiwyg = "true";
defparam \regs[30][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N31
dffeas \regs[13][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][11] .is_wysiwyg = "true";
defparam \regs[13][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N30
cycloneive_lcell_comb \Mux20~17 (
// Equation(s):
// \Mux20~17_combout  = (dcifimemload_21 & (((\regs[13][11]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][11]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][11]~q ),
	.datac(\regs[13][11]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux20~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~17 .lut_mask = 16'hAAE4;
defparam \Mux20~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y43_N31
dffeas \regs[22][10] (
	.clk(CLK),
	.d(\regs[22][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][10] .is_wysiwyg = "true";
defparam \regs[22][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y43_N15
dffeas \regs[26][10] (
	.clk(CLK),
	.d(\regs[26][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][10] .is_wysiwyg = "true";
defparam \regs[26][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N20
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (dcifimemload_23 & ((\regs[22][10]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[18][10]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[22][10]~q ),
	.datac(\regs[18][10]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hAAD8;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N30
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (dcifimemload_24 & ((\Mux21~2_combout  & ((\regs[30][10]~q ))) # (!\Mux21~2_combout  & (\regs[26][10]~q )))) # (!dcifimemload_24 & (((\Mux21~2_combout ))))

	.dataa(\regs[26][10]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[30][10]~q ),
	.datad(\Mux21~2_combout ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hF388;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y45_N23
dffeas \regs[28][9] (
	.clk(CLK),
	.d(\regs[28][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][9] .is_wysiwyg = "true";
defparam \regs[28][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N12
cycloneive_lcell_comb \Mux22~10 (
// Equation(s):
// \Mux22~10_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\regs[10][9]~q )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\regs[8][9]~q ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[10][9]~q ),
	.datad(\regs[8][9]~q ),
	.cin(gnd),
	.combout(\Mux22~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~10 .lut_mask = 16'hB9A8;
defparam \Mux22~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N27
dffeas \regs[26][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][8] .is_wysiwyg = "true";
defparam \regs[26][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N26
cycloneive_lcell_comb \Mux55~2 (
// Equation(s):
// \Mux55~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[26][8]~q ))) # (!dcifimemload_19 & (\regs[18][8]~q ))))

	.dataa(\regs[18][8]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[26][8]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux55~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~2 .lut_mask = 16'hFC22;
defparam \Mux55~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N13
dffeas \regs[23][8] (
	.clk(CLK),
	.d(\regs[23][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][8] .is_wysiwyg = "true";
defparam \regs[23][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N30
cycloneive_lcell_comb \Mux56~2 (
// Equation(s):
// \Mux56~2_combout  = (dcifimemload_18 & (((\regs[22][7]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[18][7]~q  & ((!dcifimemload_19))))

	.dataa(\regs[18][7]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[22][7]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~2 .lut_mask = 16'hCCE2;
defparam \Mux56~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N23
dffeas \regs[26][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][6] .is_wysiwyg = "true";
defparam \regs[26][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N22
cycloneive_lcell_comb \Mux57~2 (
// Equation(s):
// \Mux57~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[26][6]~q ))) # (!dcifimemload_19 & (\regs[18][6]~q ))))

	.dataa(\regs[18][6]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[26][6]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~2 .lut_mask = 16'hFC22;
defparam \Mux57~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N7
dffeas \regs[8][6] (
	.clk(CLK),
	.d(\regs[8][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][6] .is_wysiwyg = "true";
defparam \regs[8][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N13
dffeas \regs[17][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][5] .is_wysiwyg = "true";
defparam \regs[17][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N11
dffeas \regs[18][5] (
	.clk(CLK),
	.d(\regs[18][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][5] .is_wysiwyg = "true";
defparam \regs[18][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N7
dffeas \regs[30][5] (
	.clk(CLK),
	.d(\regs[30][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][5] .is_wysiwyg = "true";
defparam \regs[30][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N7
dffeas \regs[19][5] (
	.clk(CLK),
	.d(\regs[19][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][5] .is_wysiwyg = "true";
defparam \regs[19][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N30
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[21][5]~q )) # (!dcifimemload_23 & ((\regs[17][5]~q )))))

	.dataa(\regs[21][5]~q ),
	.datab(\regs[17][5]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hFA0C;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N22
cycloneive_lcell_comb \Mux26~7 (
// Equation(s):
// \Mux26~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[23][5]~q )) # (!dcifimemload_23 & ((\regs[19][5]~q )))))

	.dataa(\regs[23][5]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[19][5]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~7 .lut_mask = 16'hEE30;
defparam \Mux26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y41_N23
dffeas \regs[24][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][4] .is_wysiwyg = "true";
defparam \regs[24][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N9
dffeas \regs[16][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][4] .is_wysiwyg = "true";
defparam \regs[16][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N22
cycloneive_lcell_comb \Mux59~4 (
// Equation(s):
// \Mux59~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[24][4]~q ))) # (!dcifimemload_19 & (\regs[16][4]~q ))))

	.dataa(\regs[16][4]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[24][4]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux59~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~4 .lut_mask = 16'hFC22;
defparam \Mux59~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N26
cycloneive_lcell_comb \Mux59~12 (
// Equation(s):
// \Mux59~12_combout  = (dcifimemload_16 & (((\regs[5][4]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][4]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][4]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[5][4]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux59~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~12 .lut_mask = 16'hCCE2;
defparam \Mux59~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N8
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (dcifimemload_23 & ((\regs[20][4]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[16][4]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[20][4]~q ),
	.datac(\regs[16][4]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'hAAD8;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N30
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (dcifimemload_24 & ((\Mux27~4_combout  & ((\regs[28][4]~q ))) # (!\Mux27~4_combout  & (\regs[24][4]~q )))) # (!dcifimemload_24 & (((\Mux27~4_combout ))))

	.dataa(\regs[24][4]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[28][4]~q ),
	.datad(\Mux27~4_combout ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hF388;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N30
cycloneive_lcell_comb \Mux27~14 (
// Equation(s):
// \Mux27~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][4]~q ))) # (!dcifimemload_22 & (\regs[1][4]~q ))))

	.dataa(\regs[1][4]~q ),
	.datab(\regs[3][4]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux27~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~14 .lut_mask = 16'hC0A0;
defparam \Mux27~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N26
cycloneive_lcell_comb \Mux27~15 (
// Equation(s):
// \Mux27~15_combout  = (\Mux27~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][4]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[2][4]~q ),
	.datad(\Mux27~14_combout ),
	.cin(gnd),
	.combout(\Mux27~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~15 .lut_mask = 16'hFF20;
defparam \Mux27~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N26
cycloneive_lcell_comb \Mux60~4 (
// Equation(s):
// \Mux60~4_combout  = (dcifimemload_18 & (((\regs[20][3]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[16][3]~q  & ((!dcifimemload_19))))

	.dataa(\regs[16][3]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[20][3]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux60~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~4 .lut_mask = 16'hCCE2;
defparam \Mux60~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N25
dffeas \regs[27][3] (
	.clk(CLK),
	.d(\regs[27][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][3] .is_wysiwyg = "true";
defparam \regs[27][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N2
cycloneive_lcell_comb \Mux28~14 (
// Equation(s):
// \Mux28~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\regs[3][3]~q )) # (!dcifimemload_22 & ((\regs[1][3]~q )))))

	.dataa(\regs[3][3]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[1][3]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux28~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~14 .lut_mask = 16'h88C0;
defparam \Mux28~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N6
cycloneive_lcell_comb \Mux28~15 (
// Equation(s):
// \Mux28~15_combout  = (\Mux28~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][3]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[2][3]~q ),
	.datad(\Mux28~14_combout ),
	.cin(gnd),
	.combout(\Mux28~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~15 .lut_mask = 16'hFF20;
defparam \Mux28~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N27
dffeas \regs[4][31] (
	.clk(CLK),
	.d(\regs[4][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][31] .is_wysiwyg = "true";
defparam \regs[4][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y41_N11
dffeas \regs[25][31] (
	.clk(CLK),
	.d(\regs[25][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][31] .is_wysiwyg = "true";
defparam \regs[25][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N7
dffeas \regs[27][31] (
	.clk(CLK),
	.d(\regs[27][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][31] .is_wysiwyg = "true";
defparam \regs[27][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N22
cycloneive_lcell_comb \regs~12 (
// Equation(s):
// \regs~12_combout  = (cuifRegSel_0) # ((\regs~11_combout  & (\Add1~50_combout )) # (!\regs~11_combout  & ((Selector0))))

	.dataa(Add117),
	.datab(cuifRegSel_0),
	.datac(\regs~11_combout ),
	.datad(Selector0),
	.cin(gnd),
	.combout(\regs~12_combout ),
	.cout());
// synopsys translate_off
defparam \regs~12 .lut_mask = 16'hEFEC;
defparam \regs~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N30
cycloneive_lcell_comb \regs~15 (
// Equation(s):
// \regs~15_combout  = (cuifRegSel_11) # ((\regs~14_combout  & (ramiframload_261)) # (!\regs~14_combout  & ((Selector0))))

	.dataa(ramiframload_26),
	.datab(Selector0),
	.datac(cuifRegSel_11),
	.datad(\regs~14_combout ),
	.cin(gnd),
	.combout(\regs~15_combout ),
	.cout());
// synopsys translate_off
defparam \regs~15 .lut_mask = 16'hFAFC;
defparam \regs~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N30
cycloneive_lcell_comb \regs~59 (
// Equation(s):
// \regs~59_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_3)) # (!cuifRegSel_0 & ((Mux281)))))

	.dataa(ramiframload_3),
	.datab(cuifRegSel_11),
	.datac(Mux281),
	.datad(cuifRegSel_0),
	.cin(gnd),
	.combout(\regs~59_combout ),
	.cout());
// synopsys translate_off
defparam \regs~59 .lut_mask = 16'h2230;
defparam \regs~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N12
cycloneive_lcell_comb \regs[21][0]~feeder (
// Equation(s):
// \regs[21][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~5_combout ),
	.cin(gnd),
	.combout(\regs[21][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][0]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N26
cycloneive_lcell_comb \regs[26][1]~feeder (
// Equation(s):
// \regs[26][1]~feeder_combout  = \regs~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[26][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][1]~feeder .lut_mask = 16'hF0F0;
defparam \regs[26][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N10
cycloneive_lcell_comb \regs[27][1]~feeder (
// Equation(s):
// \regs[27][1]~feeder_combout  = \regs~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][1]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N24
cycloneive_lcell_comb \regs[18][30]~feeder (
// Equation(s):
// \regs[18][30]~feeder_combout  = \regs~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[18][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[18][30]~feeder .lut_mask = 16'hF0F0;
defparam \regs[18][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N22
cycloneive_lcell_comb \regs[17][30]~feeder (
// Equation(s):
// \regs[17][30]~feeder_combout  = \regs~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[17][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][30]~feeder .lut_mask = 16'hF0F0;
defparam \regs[17][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N30
cycloneive_lcell_comb \regs[26][29]~feeder (
// Equation(s):
// \regs[26][29]~feeder_combout  = \regs~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[26][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][29]~feeder .lut_mask = 16'hF0F0;
defparam \regs[26][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N22
cycloneive_lcell_comb \regs[5][24]~feeder (
// Equation(s):
// \regs[5][24]~feeder_combout  = \regs~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~22_combout ),
	.cin(gnd),
	.combout(\regs[5][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[5][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N26
cycloneive_lcell_comb \regs[8][19]~feeder (
// Equation(s):
// \regs[8][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~27_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[8][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[8][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N12
cycloneive_lcell_comb \regs[11][17]~feeder (
// Equation(s):
// \regs[11][17]~feeder_combout  = \regs~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~29_combout ),
	.cin(gnd),
	.combout(\regs[11][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][17]~feeder .lut_mask = 16'hFF00;
defparam \regs[11][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N8
cycloneive_lcell_comb \regs[8][17]~feeder (
// Equation(s):
// \regs[8][17]~feeder_combout  = \regs~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~29_combout ),
	.cin(gnd),
	.combout(\regs[8][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][17]~feeder .lut_mask = 16'hFF00;
defparam \regs[8][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N12
cycloneive_lcell_comb \regs[17][15]~feeder (
// Equation(s):
// \regs[17][15]~feeder_combout  = \regs~32_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~32_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[17][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][15]~feeder .lut_mask = 16'hF0F0;
defparam \regs[17][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N10
cycloneive_lcell_comb \regs[22][14]~feeder (
// Equation(s):
// \regs[22][14]~feeder_combout  = \regs~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~34_combout ),
	.cin(gnd),
	.combout(\regs[22][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][14]~feeder .lut_mask = 16'hFF00;
defparam \regs[22][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N6
cycloneive_lcell_comb \regs[26][14]~feeder (
// Equation(s):
// \regs[26][14]~feeder_combout  = \regs~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~34_combout ),
	.cin(gnd),
	.combout(\regs[26][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][14]~feeder .lut_mask = 16'hFF00;
defparam \regs[26][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N22
cycloneive_lcell_comb \regs[3][13]~feeder (
// Equation(s):
// \regs[3][13]~feeder_combout  = \regs~36_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~36_combout ),
	.cin(gnd),
	.combout(\regs[3][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N6
cycloneive_lcell_comb \regs[24][12]~feeder (
// Equation(s):
// \regs[24][12]~feeder_combout  = \regs~38_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~38_combout ),
	.cin(gnd),
	.combout(\regs[24][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][12]~feeder .lut_mask = 16'hFF00;
defparam \regs[24][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N30
cycloneive_lcell_comb \regs[30][11]~feeder (
// Equation(s):
// \regs[30][11]~feeder_combout  = \regs~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~40_combout ),
	.cin(gnd),
	.combout(\regs[30][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[30][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[30][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N30
cycloneive_lcell_comb \regs[22][10]~feeder (
// Equation(s):
// \regs[22][10]~feeder_combout  = \regs~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~42_combout ),
	.cin(gnd),
	.combout(\regs[22][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][10]~feeder .lut_mask = 16'hFF00;
defparam \regs[22][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N14
cycloneive_lcell_comb \regs[26][10]~feeder (
// Equation(s):
// \regs[26][10]~feeder_combout  = \regs~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~42_combout ),
	.cin(gnd),
	.combout(\regs[26][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][10]~feeder .lut_mask = 16'hFF00;
defparam \regs[26][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N22
cycloneive_lcell_comb \regs[28][9]~feeder (
// Equation(s):
// \regs[28][9]~feeder_combout  = \regs~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[28][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][9]~feeder .lut_mask = 16'hF0F0;
defparam \regs[28][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N12
cycloneive_lcell_comb \regs[23][8]~feeder (
// Equation(s):
// \regs[23][8]~feeder_combout  = \regs~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~46_combout ),
	.cin(gnd),
	.combout(\regs[23][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][8]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N6
cycloneive_lcell_comb \regs[8][6]~feeder (
// Equation(s):
// \regs[8][6]~feeder_combout  = \regs~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[8][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[8][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N6
cycloneive_lcell_comb \regs[19][5]~feeder (
// Equation(s):
// \regs[19][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[19][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[19][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N10
cycloneive_lcell_comb \regs[18][5]~feeder (
// Equation(s):
// \regs[18][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[18][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[18][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[18][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N6
cycloneive_lcell_comb \regs[30][5]~feeder (
// Equation(s):
// \regs[30][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[30][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[30][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[30][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N24
cycloneive_lcell_comb \regs[27][3]~feeder (
// Equation(s):
// \regs[27][3]~feeder_combout  = \regs~60_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~60_combout ),
	.cin(gnd),
	.combout(\regs[27][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][3]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N10
cycloneive_lcell_comb \regs[25][31]~feeder (
// Equation(s):
// \regs[25][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~63_combout ),
	.cin(gnd),
	.combout(\regs[25][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[25][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[25][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N6
cycloneive_lcell_comb \regs[27][31]~feeder (
// Equation(s):
// \regs[27][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~63_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][31]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N26
cycloneive_lcell_comb \regs[4][31]~feeder (
// Equation(s):
// \regs[4][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~63_combout ),
	.cin(gnd),
	.combout(\regs[4][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[4][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[4][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N0
cycloneive_lcell_comb \Mux63~9 (
// Equation(s):
// Mux63 = (\Mux63~6_combout  & (((\Mux63~8_combout ) # (!dcifimemload_16)))) # (!\Mux63~6_combout  & (\Mux63~1_combout  & (dcifimemload_16)))

	.dataa(\Mux63~6_combout ),
	.datab(\Mux63~1_combout ),
	.datac(dcifimemload_16),
	.datad(\Mux63~8_combout ),
	.cin(gnd),
	.combout(Mux63),
	.cout());
// synopsys translate_off
defparam \Mux63~9 .lut_mask = 16'hEA4A;
defparam \Mux63~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N24
cycloneive_lcell_comb \Mux63~19 (
// Equation(s):
// Mux631 = (dcifimemload_19 & ((\Mux63~16_combout  & ((\Mux63~18_combout ))) # (!\Mux63~16_combout  & (\Mux63~11_combout )))) # (!dcifimemload_19 & (((\Mux63~16_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux63~11_combout ),
	.datac(\Mux63~18_combout ),
	.datad(\Mux63~16_combout ),
	.cin(gnd),
	.combout(Mux631),
	.cout());
// synopsys translate_off
defparam \Mux63~19 .lut_mask = 16'hF588;
defparam \Mux63~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N0
cycloneive_lcell_comb \Mux30~20 (
// Equation(s):
// Mux30 = (dcifimemload_25 & (\Mux30~9_combout )) # (!dcifimemload_25 & ((\Mux30~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux30~9_combout ),
	.datad(\Mux30~19_combout ),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~20 .lut_mask = 16'hF5A0;
defparam \Mux30~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N18
cycloneive_lcell_comb \Mux33~9 (
// Equation(s):
// Mux33 = (dcifimemload_16 & ((\Mux33~6_combout  & (\Mux33~8_combout )) # (!\Mux33~6_combout  & ((\Mux33~1_combout ))))) # (!dcifimemload_16 & (((\Mux33~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux33~8_combout ),
	.datac(\Mux33~1_combout ),
	.datad(\Mux33~6_combout ),
	.cin(gnd),
	.combout(Mux33),
	.cout());
// synopsys translate_off
defparam \Mux33~9 .lut_mask = 16'hDDA0;
defparam \Mux33~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N22
cycloneive_lcell_comb \Mux33~19 (
// Equation(s):
// Mux331 = (dcifimemload_19 & ((\Mux33~16_combout  & (\Mux33~18_combout )) # (!\Mux33~16_combout  & ((\Mux33~11_combout ))))) # (!dcifimemload_19 & (((\Mux33~16_combout ))))

	.dataa(\Mux33~18_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux33~11_combout ),
	.datad(\Mux33~16_combout ),
	.cin(gnd),
	.combout(Mux331),
	.cout());
// synopsys translate_off
defparam \Mux33~19 .lut_mask = 16'hBBC0;
defparam \Mux33~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N22
cycloneive_lcell_comb \Mux1~20 (
// Equation(s):
// Mux1 = (dcifimemload_25 & ((\Mux1~9_combout ))) # (!dcifimemload_25 & (\Mux1~19_combout ))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux1~19_combout ),
	.datad(\Mux1~9_combout ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~20 .lut_mask = 16'hFA50;
defparam \Mux1~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N16
cycloneive_lcell_comb \Mux34~9 (
// Equation(s):
// Mux34 = (dcifimemload_16 & ((\Mux34~6_combout  & (\Mux34~8_combout )) # (!\Mux34~6_combout  & ((\Mux34~1_combout ))))) # (!dcifimemload_16 & (((\Mux34~6_combout ))))

	.dataa(\Mux34~8_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux34~1_combout ),
	.datad(\Mux34~6_combout ),
	.cin(gnd),
	.combout(Mux34),
	.cout());
// synopsys translate_off
defparam \Mux34~9 .lut_mask = 16'hBBC0;
defparam \Mux34~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N20
cycloneive_lcell_comb \Mux34~19 (
// Equation(s):
// Mux341 = (dcifimemload_18 & ((\Mux34~16_combout  & ((\Mux34~18_combout ))) # (!\Mux34~16_combout  & (\Mux34~11_combout )))) # (!dcifimemload_18 & (((\Mux34~16_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux34~11_combout ),
	.datac(\Mux34~18_combout ),
	.datad(\Mux34~16_combout ),
	.cin(gnd),
	.combout(Mux341),
	.cout());
// synopsys translate_off
defparam \Mux34~19 .lut_mask = 16'hF588;
defparam \Mux34~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N2
cycloneive_lcell_comb \Mux2~20 (
// Equation(s):
// Mux2 = (dcifimemload_25 & (\Mux2~9_combout )) # (!dcifimemload_25 & ((\Mux2~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux2~9_combout ),
	.datad(\Mux2~19_combout ),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~20 .lut_mask = 16'hF5A0;
defparam \Mux2~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N0
cycloneive_lcell_comb \Mux35~9 (
// Equation(s):
// Mux35 = (\Mux35~6_combout  & (((\Mux35~8_combout )) # (!dcifimemload_16))) # (!\Mux35~6_combout  & (dcifimemload_16 & ((\Mux35~1_combout ))))

	.dataa(\Mux35~6_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux35~8_combout ),
	.datad(\Mux35~1_combout ),
	.cin(gnd),
	.combout(Mux35),
	.cout());
// synopsys translate_off
defparam \Mux35~9 .lut_mask = 16'hE6A2;
defparam \Mux35~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N6
cycloneive_lcell_comb \Mux35~19 (
// Equation(s):
// Mux351 = (dcifimemload_19 & ((\Mux35~16_combout  & (\Mux35~18_combout )) # (!\Mux35~16_combout  & ((\Mux35~11_combout ))))) # (!dcifimemload_19 & (((\Mux35~16_combout ))))

	.dataa(\Mux35~18_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux35~11_combout ),
	.datad(\Mux35~16_combout ),
	.cin(gnd),
	.combout(Mux351),
	.cout());
// synopsys translate_off
defparam \Mux35~19 .lut_mask = 16'hBBC0;
defparam \Mux35~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N6
cycloneive_lcell_comb \Mux3~20 (
// Equation(s):
// Mux3 = (dcifimemload_25 & ((\Mux3~9_combout ))) # (!dcifimemload_25 & (\Mux3~19_combout ))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux3~19_combout ),
	.datad(\Mux3~9_combout ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~20 .lut_mask = 16'hFC30;
defparam \Mux3~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N24
cycloneive_lcell_comb \Mux36~9 (
// Equation(s):
// Mux36 = (\Mux36~6_combout  & (((\Mux36~8_combout )) # (!dcifimemload_16))) # (!\Mux36~6_combout  & (dcifimemload_16 & ((\Mux36~1_combout ))))

	.dataa(\Mux36~6_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux36~8_combout ),
	.datad(\Mux36~1_combout ),
	.cin(gnd),
	.combout(Mux36),
	.cout());
// synopsys translate_off
defparam \Mux36~9 .lut_mask = 16'hE6A2;
defparam \Mux36~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N12
cycloneive_lcell_comb \Mux36~19 (
// Equation(s):
// Mux361 = (dcifimemload_18 & ((\Mux36~16_combout  & ((\Mux36~18_combout ))) # (!\Mux36~16_combout  & (\Mux36~11_combout )))) # (!dcifimemload_18 & (((\Mux36~16_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux36~11_combout ),
	.datac(\Mux36~16_combout ),
	.datad(\Mux36~18_combout ),
	.cin(gnd),
	.combout(Mux361),
	.cout());
// synopsys translate_off
defparam \Mux36~19 .lut_mask = 16'hF858;
defparam \Mux36~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N2
cycloneive_lcell_comb \Mux4~20 (
// Equation(s):
// Mux4 = (dcifimemload_25 & (\Mux4~9_combout )) # (!dcifimemload_25 & ((\Mux4~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux4~9_combout ),
	.datad(\Mux4~19_combout ),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~20 .lut_mask = 16'hF3C0;
defparam \Mux4~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N10
cycloneive_lcell_comb \Mux37~9 (
// Equation(s):
// Mux37 = (dcifimemload_16 & ((\Mux37~6_combout  & (\Mux37~8_combout )) # (!\Mux37~6_combout  & ((\Mux37~1_combout ))))) # (!dcifimemload_16 & (\Mux37~6_combout ))

	.dataa(dcifimemload_16),
	.datab(\Mux37~6_combout ),
	.datac(\Mux37~8_combout ),
	.datad(\Mux37~1_combout ),
	.cin(gnd),
	.combout(Mux37),
	.cout());
// synopsys translate_off
defparam \Mux37~9 .lut_mask = 16'hE6C4;
defparam \Mux37~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N4
cycloneive_lcell_comb \Mux37~19 (
// Equation(s):
// Mux371 = (dcifimemload_19 & ((\Mux37~16_combout  & ((\Mux37~18_combout ))) # (!\Mux37~16_combout  & (\Mux37~11_combout )))) # (!dcifimemload_19 & (((\Mux37~16_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux37~11_combout ),
	.datac(\Mux37~18_combout ),
	.datad(\Mux37~16_combout ),
	.cin(gnd),
	.combout(Mux371),
	.cout());
// synopsys translate_off
defparam \Mux37~19 .lut_mask = 16'hF588;
defparam \Mux37~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N10
cycloneive_lcell_comb \Mux5~20 (
// Equation(s):
// Mux5 = (dcifimemload_25 & (\Mux5~9_combout )) # (!dcifimemload_25 & ((\Mux5~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux5~9_combout ),
	.datad(\Mux5~19_combout ),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~20 .lut_mask = 16'hF5A0;
defparam \Mux5~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N18
cycloneive_lcell_comb \Mux38~9 (
// Equation(s):
// Mux38 = (\Mux38~6_combout  & (((\Mux38~8_combout )) # (!dcifimemload_16))) # (!\Mux38~6_combout  & (dcifimemload_16 & (\Mux38~1_combout )))

	.dataa(\Mux38~6_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux38~1_combout ),
	.datad(\Mux38~8_combout ),
	.cin(gnd),
	.combout(Mux38),
	.cout());
// synopsys translate_off
defparam \Mux38~9 .lut_mask = 16'hEA62;
defparam \Mux38~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N30
cycloneive_lcell_comb \Mux38~19 (
// Equation(s):
// Mux381 = (dcifimemload_18 & ((\Mux38~16_combout  & ((\Mux38~18_combout ))) # (!\Mux38~16_combout  & (\Mux38~11_combout )))) # (!dcifimemload_18 & (((\Mux38~16_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux38~11_combout ),
	.datac(\Mux38~18_combout ),
	.datad(\Mux38~16_combout ),
	.cin(gnd),
	.combout(Mux381),
	.cout());
// synopsys translate_off
defparam \Mux38~19 .lut_mask = 16'hF588;
defparam \Mux38~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N22
cycloneive_lcell_comb \Mux6~20 (
// Equation(s):
// Mux6 = (dcifimemload_25 & (\Mux6~9_combout )) # (!dcifimemload_25 & ((\Mux6~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux6~9_combout ),
	.datad(\Mux6~19_combout ),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~20 .lut_mask = 16'hF5A0;
defparam \Mux6~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N18
cycloneive_lcell_comb \Mux39~9 (
// Equation(s):
// Mux39 = (dcifimemload_16 & ((\Mux39~6_combout  & (\Mux39~8_combout )) # (!\Mux39~6_combout  & ((\Mux39~1_combout ))))) # (!dcifimemload_16 & (((\Mux39~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux39~8_combout ),
	.datac(\Mux39~1_combout ),
	.datad(\Mux39~6_combout ),
	.cin(gnd),
	.combout(Mux39),
	.cout());
// synopsys translate_off
defparam \Mux39~9 .lut_mask = 16'hDDA0;
defparam \Mux39~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N30
cycloneive_lcell_comb \Mux39~19 (
// Equation(s):
// Mux391 = (dcifimemload_19 & ((\Mux39~16_combout  & (\Mux39~18_combout )) # (!\Mux39~16_combout  & ((\Mux39~11_combout ))))) # (!dcifimemload_19 & (((\Mux39~16_combout ))))

	.dataa(\Mux39~18_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux39~11_combout ),
	.datad(\Mux39~16_combout ),
	.cin(gnd),
	.combout(Mux391),
	.cout());
// synopsys translate_off
defparam \Mux39~19 .lut_mask = 16'hBBC0;
defparam \Mux39~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N10
cycloneive_lcell_comb \Mux7~20 (
// Equation(s):
// Mux7 = (dcifimemload_25 & (\Mux7~9_combout )) # (!dcifimemload_25 & ((\Mux7~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux7~9_combout ),
	.datad(\Mux7~19_combout ),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~20 .lut_mask = 16'hF3C0;
defparam \Mux7~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N22
cycloneive_lcell_comb \Mux40~9 (
// Equation(s):
// Mux40 = (dcifimemload_16 & ((\Mux40~6_combout  & ((\Mux40~8_combout ))) # (!\Mux40~6_combout  & (\Mux40~1_combout )))) # (!dcifimemload_16 & (((\Mux40~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux40~1_combout ),
	.datac(\Mux40~6_combout ),
	.datad(\Mux40~8_combout ),
	.cin(gnd),
	.combout(Mux40),
	.cout());
// synopsys translate_off
defparam \Mux40~9 .lut_mask = 16'hF858;
defparam \Mux40~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N26
cycloneive_lcell_comb \Mux40~19 (
// Equation(s):
// Mux401 = (dcifimemload_18 & ((\Mux40~16_combout  & ((\Mux40~18_combout ))) # (!\Mux40~16_combout  & (\Mux40~11_combout )))) # (!dcifimemload_18 & (((\Mux40~16_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux40~11_combout ),
	.datac(\Mux40~18_combout ),
	.datad(\Mux40~16_combout ),
	.cin(gnd),
	.combout(Mux401),
	.cout());
// synopsys translate_off
defparam \Mux40~19 .lut_mask = 16'hF588;
defparam \Mux40~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N14
cycloneive_lcell_comb \Mux8~20 (
// Equation(s):
// Mux8 = (dcifimemload_25 & (\Mux8~9_combout )) # (!dcifimemload_25 & ((\Mux8~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux8~9_combout ),
	.datad(\Mux8~19_combout ),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~20 .lut_mask = 16'hF3C0;
defparam \Mux8~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N6
cycloneive_lcell_comb \Mux41~9 (
// Equation(s):
// Mux41 = (dcifimemload_16 & ((\Mux41~6_combout  & ((\Mux41~8_combout ))) # (!\Mux41~6_combout  & (\Mux41~1_combout )))) # (!dcifimemload_16 & (((\Mux41~6_combout ))))

	.dataa(\Mux41~1_combout ),
	.datab(\Mux41~8_combout ),
	.datac(dcifimemload_16),
	.datad(\Mux41~6_combout ),
	.cin(gnd),
	.combout(Mux41),
	.cout());
// synopsys translate_off
defparam \Mux41~9 .lut_mask = 16'hCFA0;
defparam \Mux41~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N18
cycloneive_lcell_comb \Mux41~19 (
// Equation(s):
// Mux411 = (dcifimemload_19 & ((\Mux41~16_combout  & ((\Mux41~18_combout ))) # (!\Mux41~16_combout  & (\Mux41~11_combout )))) # (!dcifimemload_19 & (((\Mux41~16_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux41~11_combout ),
	.datac(\Mux41~16_combout ),
	.datad(\Mux41~18_combout ),
	.cin(gnd),
	.combout(Mux411),
	.cout());
// synopsys translate_off
defparam \Mux41~19 .lut_mask = 16'hF858;
defparam \Mux41~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N28
cycloneive_lcell_comb \Mux9~20 (
// Equation(s):
// Mux9 = (dcifimemload_25 & (\Mux9~9_combout )) # (!dcifimemload_25 & ((\Mux9~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux9~9_combout ),
	.datad(\Mux9~19_combout ),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~20 .lut_mask = 16'hF5A0;
defparam \Mux9~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N24
cycloneive_lcell_comb \Mux42~9 (
// Equation(s):
// Mux42 = (dcifimemload_16 & ((\Mux42~6_combout  & (\Mux42~8_combout )) # (!\Mux42~6_combout  & ((\Mux42~1_combout ))))) # (!dcifimemload_16 & (((\Mux42~6_combout ))))

	.dataa(\Mux42~8_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux42~1_combout ),
	.datad(\Mux42~6_combout ),
	.cin(gnd),
	.combout(Mux42),
	.cout());
// synopsys translate_off
defparam \Mux42~9 .lut_mask = 16'hBBC0;
defparam \Mux42~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N8
cycloneive_lcell_comb \Mux42~19 (
// Equation(s):
// Mux421 = (\Mux42~16_combout  & (((\Mux42~18_combout )) # (!dcifimemload_18))) # (!\Mux42~16_combout  & (dcifimemload_18 & (\Mux42~11_combout )))

	.dataa(\Mux42~16_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux42~11_combout ),
	.datad(\Mux42~18_combout ),
	.cin(gnd),
	.combout(Mux421),
	.cout());
// synopsys translate_off
defparam \Mux42~19 .lut_mask = 16'hEA62;
defparam \Mux42~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N28
cycloneive_lcell_comb \Mux10~20 (
// Equation(s):
// Mux10 = (dcifimemload_25 & (\Mux10~9_combout )) # (!dcifimemload_25 & ((\Mux10~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux10~9_combout ),
	.datad(\Mux10~19_combout ),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~20 .lut_mask = 16'hF5A0;
defparam \Mux10~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N10
cycloneive_lcell_comb \Mux43~9 (
// Equation(s):
// Mux43 = (dcifimemload_16 & ((\Mux43~6_combout  & (\Mux43~8_combout )) # (!\Mux43~6_combout  & ((\Mux43~1_combout ))))) # (!dcifimemload_16 & (((\Mux43~6_combout ))))

	.dataa(\Mux43~8_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux43~6_combout ),
	.datad(\Mux43~1_combout ),
	.cin(gnd),
	.combout(Mux43),
	.cout());
// synopsys translate_off
defparam \Mux43~9 .lut_mask = 16'hBCB0;
defparam \Mux43~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N28
cycloneive_lcell_comb \Mux43~19 (
// Equation(s):
// Mux431 = (dcifimemload_19 & ((\Mux43~16_combout  & (\Mux43~18_combout )) # (!\Mux43~16_combout  & ((\Mux43~11_combout ))))) # (!dcifimemload_19 & (((\Mux43~16_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux43~18_combout ),
	.datac(\Mux43~11_combout ),
	.datad(\Mux43~16_combout ),
	.cin(gnd),
	.combout(Mux431),
	.cout());
// synopsys translate_off
defparam \Mux43~19 .lut_mask = 16'hDDA0;
defparam \Mux43~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N18
cycloneive_lcell_comb \Mux11~20 (
// Equation(s):
// Mux11 = (dcifimemload_25 & (\Mux11~9_combout )) # (!dcifimemload_25 & ((\Mux11~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux11~9_combout ),
	.datad(\Mux11~19_combout ),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux11~20 .lut_mask = 16'hF5A0;
defparam \Mux11~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N2
cycloneive_lcell_comb \Mux44~9 (
// Equation(s):
// Mux44 = (dcifimemload_16 & ((\Mux44~6_combout  & (\Mux44~8_combout )) # (!\Mux44~6_combout  & ((\Mux44~1_combout ))))) # (!dcifimemload_16 & (((\Mux44~6_combout ))))

	.dataa(\Mux44~8_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux44~6_combout ),
	.datad(\Mux44~1_combout ),
	.cin(gnd),
	.combout(Mux44),
	.cout());
// synopsys translate_off
defparam \Mux44~9 .lut_mask = 16'hBCB0;
defparam \Mux44~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N0
cycloneive_lcell_comb \Mux44~19 (
// Equation(s):
// Mux441 = (dcifimemload_18 & ((\Mux44~16_combout  & (\Mux44~18_combout )) # (!\Mux44~16_combout  & ((\Mux44~11_combout ))))) # (!dcifimemload_18 & (((\Mux44~16_combout ))))

	.dataa(\Mux44~18_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux44~16_combout ),
	.datad(\Mux44~11_combout ),
	.cin(gnd),
	.combout(Mux441),
	.cout());
// synopsys translate_off
defparam \Mux44~19 .lut_mask = 16'hBCB0;
defparam \Mux44~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N2
cycloneive_lcell_comb \Mux12~20 (
// Equation(s):
// Mux12 = (dcifimemload_25 & (\Mux12~9_combout )) # (!dcifimemload_25 & ((\Mux12~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux12~9_combout ),
	.datad(\Mux12~19_combout ),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~20 .lut_mask = 16'hF5A0;
defparam \Mux12~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N10
cycloneive_lcell_comb \Mux45~9 (
// Equation(s):
// Mux45 = (dcifimemload_16 & ((\Mux45~6_combout  & (\Mux45~8_combout )) # (!\Mux45~6_combout  & ((\Mux45~1_combout ))))) # (!dcifimemload_16 & (\Mux45~6_combout ))

	.dataa(dcifimemload_16),
	.datab(\Mux45~6_combout ),
	.datac(\Mux45~8_combout ),
	.datad(\Mux45~1_combout ),
	.cin(gnd),
	.combout(Mux45),
	.cout());
// synopsys translate_off
defparam \Mux45~9 .lut_mask = 16'hE6C4;
defparam \Mux45~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N18
cycloneive_lcell_comb \Mux45~19 (
// Equation(s):
// Mux451 = (dcifimemload_19 & ((\Mux45~16_combout  & (\Mux45~18_combout )) # (!\Mux45~16_combout  & ((\Mux45~11_combout ))))) # (!dcifimemload_19 & (((\Mux45~16_combout ))))

	.dataa(\Mux45~18_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux45~11_combout ),
	.datad(\Mux45~16_combout ),
	.cin(gnd),
	.combout(Mux451),
	.cout());
// synopsys translate_off
defparam \Mux45~19 .lut_mask = 16'hBBC0;
defparam \Mux45~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N6
cycloneive_lcell_comb \Mux13~20 (
// Equation(s):
// Mux13 = (dcifimemload_25 & (\Mux13~9_combout )) # (!dcifimemload_25 & ((\Mux13~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux13~9_combout ),
	.datad(\Mux13~19_combout ),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~20 .lut_mask = 16'hF3C0;
defparam \Mux13~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N14
cycloneive_lcell_comb \Mux46~9 (
// Equation(s):
// Mux46 = (dcifimemload_16 & ((\Mux46~6_combout  & ((\Mux46~8_combout ))) # (!\Mux46~6_combout  & (\Mux46~1_combout )))) # (!dcifimemload_16 & (((\Mux46~6_combout ))))

	.dataa(\Mux46~1_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux46~8_combout ),
	.datad(\Mux46~6_combout ),
	.cin(gnd),
	.combout(Mux46),
	.cout());
// synopsys translate_off
defparam \Mux46~9 .lut_mask = 16'hF388;
defparam \Mux46~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N26
cycloneive_lcell_comb \Mux46~19 (
// Equation(s):
// Mux461 = (dcifimemload_18 & ((\Mux46~16_combout  & (\Mux46~18_combout )) # (!\Mux46~16_combout  & ((\Mux46~11_combout ))))) # (!dcifimemload_18 & (((\Mux46~16_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux46~18_combout ),
	.datac(\Mux46~11_combout ),
	.datad(\Mux46~16_combout ),
	.cin(gnd),
	.combout(Mux461),
	.cout());
// synopsys translate_off
defparam \Mux46~19 .lut_mask = 16'hDDA0;
defparam \Mux46~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N2
cycloneive_lcell_comb \Mux14~20 (
// Equation(s):
// Mux14 = (dcifimemload_25 & (\Mux14~9_combout )) # (!dcifimemload_25 & ((\Mux14~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux14~9_combout ),
	.datad(\Mux14~19_combout ),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~20 .lut_mask = 16'hF3C0;
defparam \Mux14~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N0
cycloneive_lcell_comb \Mux47~9 (
// Equation(s):
// Mux47 = (dcifimemload_16 & ((\Mux47~6_combout  & ((\Mux47~8_combout ))) # (!\Mux47~6_combout  & (\Mux47~1_combout )))) # (!dcifimemload_16 & (((\Mux47~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux47~1_combout ),
	.datac(\Mux47~6_combout ),
	.datad(\Mux47~8_combout ),
	.cin(gnd),
	.combout(Mux47),
	.cout());
// synopsys translate_off
defparam \Mux47~9 .lut_mask = 16'hF858;
defparam \Mux47~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N22
cycloneive_lcell_comb \Mux47~19 (
// Equation(s):
// Mux471 = (dcifimemload_19 & ((\Mux47~16_combout  & (\Mux47~18_combout )) # (!\Mux47~16_combout  & ((\Mux47~11_combout ))))) # (!dcifimemload_19 & (((\Mux47~16_combout ))))

	.dataa(\Mux47~18_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux47~11_combout ),
	.datad(\Mux47~16_combout ),
	.cin(gnd),
	.combout(Mux471),
	.cout());
// synopsys translate_off
defparam \Mux47~19 .lut_mask = 16'hBBC0;
defparam \Mux47~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N26
cycloneive_lcell_comb \Mux15~20 (
// Equation(s):
// Mux15 = (dcifimemload_25 & ((\Mux15~9_combout ))) # (!dcifimemload_25 & (\Mux15~19_combout ))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux15~19_combout ),
	.datad(\Mux15~9_combout ),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~20 .lut_mask = 16'hFA50;
defparam \Mux15~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N16
cycloneive_lcell_comb \Mux48~9 (
// Equation(s):
// Mux48 = (\Mux48~6_combout  & (((\Mux48~8_combout )) # (!dcifimemload_16))) # (!\Mux48~6_combout  & (dcifimemload_16 & (\Mux48~1_combout )))

	.dataa(\Mux48~6_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux48~1_combout ),
	.datad(\Mux48~8_combout ),
	.cin(gnd),
	.combout(Mux48),
	.cout());
// synopsys translate_off
defparam \Mux48~9 .lut_mask = 16'hEA62;
defparam \Mux48~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N4
cycloneive_lcell_comb \Mux48~19 (
// Equation(s):
// Mux481 = (dcifimemload_18 & ((\Mux48~16_combout  & ((\Mux48~18_combout ))) # (!\Mux48~16_combout  & (\Mux48~11_combout )))) # (!dcifimemload_18 & (((\Mux48~16_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux48~11_combout ),
	.datac(\Mux48~18_combout ),
	.datad(\Mux48~16_combout ),
	.cin(gnd),
	.combout(Mux481),
	.cout());
// synopsys translate_off
defparam \Mux48~19 .lut_mask = 16'hF588;
defparam \Mux48~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N14
cycloneive_lcell_comb \Mux16~20 (
// Equation(s):
// Mux16 = (dcifimemload_25 & ((\Mux16~9_combout ))) # (!dcifimemload_25 & (\Mux16~19_combout ))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux16~19_combout ),
	.datad(\Mux16~9_combout ),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~20 .lut_mask = 16'hFA50;
defparam \Mux16~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N16
cycloneive_lcell_comb \Mux49~9 (
// Equation(s):
// Mux49 = (dcifimemload_16 & ((\Mux49~6_combout  & ((\Mux49~8_combout ))) # (!\Mux49~6_combout  & (\Mux49~1_combout )))) # (!dcifimemload_16 & (((\Mux49~6_combout ))))

	.dataa(\Mux49~1_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux49~6_combout ),
	.datad(\Mux49~8_combout ),
	.cin(gnd),
	.combout(Mux49),
	.cout());
// synopsys translate_off
defparam \Mux49~9 .lut_mask = 16'hF838;
defparam \Mux49~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N4
cycloneive_lcell_comb \Mux49~19 (
// Equation(s):
// Mux491 = (dcifimemload_19 & ((\Mux49~16_combout  & ((\Mux49~18_combout ))) # (!\Mux49~16_combout  & (\Mux49~11_combout )))) # (!dcifimemload_19 & (((\Mux49~16_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux49~11_combout ),
	.datac(\Mux49~18_combout ),
	.datad(\Mux49~16_combout ),
	.cin(gnd),
	.combout(Mux491),
	.cout());
// synopsys translate_off
defparam \Mux49~19 .lut_mask = 16'hF588;
defparam \Mux49~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N6
cycloneive_lcell_comb \Mux17~20 (
// Equation(s):
// Mux17 = (dcifimemload_25 & (\Mux17~9_combout )) # (!dcifimemload_25 & ((\Mux17~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux17~9_combout ),
	.datad(\Mux17~19_combout ),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~20 .lut_mask = 16'hF3C0;
defparam \Mux17~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N2
cycloneive_lcell_comb \Mux50~9 (
// Equation(s):
// Mux50 = (dcifimemload_16 & ((\Mux50~6_combout  & (\Mux50~8_combout )) # (!\Mux50~6_combout  & ((\Mux50~1_combout ))))) # (!dcifimemload_16 & (((\Mux50~6_combout ))))

	.dataa(\Mux50~8_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux50~6_combout ),
	.datad(\Mux50~1_combout ),
	.cin(gnd),
	.combout(Mux50),
	.cout());
// synopsys translate_off
defparam \Mux50~9 .lut_mask = 16'hBCB0;
defparam \Mux50~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N26
cycloneive_lcell_comb \Mux50~19 (
// Equation(s):
// Mux501 = (dcifimemload_18 & ((\Mux50~16_combout  & (\Mux50~18_combout )) # (!\Mux50~16_combout  & ((\Mux50~11_combout ))))) # (!dcifimemload_18 & (((\Mux50~16_combout ))))

	.dataa(\Mux50~18_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux50~11_combout ),
	.datad(\Mux50~16_combout ),
	.cin(gnd),
	.combout(Mux501),
	.cout());
// synopsys translate_off
defparam \Mux50~19 .lut_mask = 16'hBBC0;
defparam \Mux50~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N6
cycloneive_lcell_comb \Mux18~20 (
// Equation(s):
// Mux18 = (dcifimemload_25 & (\Mux18~9_combout )) # (!dcifimemload_25 & ((\Mux18~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux18~9_combout ),
	.datad(\Mux18~19_combout ),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~20 .lut_mask = 16'hF5A0;
defparam \Mux18~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N22
cycloneive_lcell_comb \Mux51~9 (
// Equation(s):
// Mux51 = (dcifimemload_16 & ((\Mux51~6_combout  & (\Mux51~8_combout )) # (!\Mux51~6_combout  & ((\Mux51~1_combout ))))) # (!dcifimemload_16 & (((\Mux51~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux51~8_combout ),
	.datac(\Mux51~1_combout ),
	.datad(\Mux51~6_combout ),
	.cin(gnd),
	.combout(Mux51),
	.cout());
// synopsys translate_off
defparam \Mux51~9 .lut_mask = 16'hDDA0;
defparam \Mux51~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N0
cycloneive_lcell_comb \Mux51~19 (
// Equation(s):
// Mux511 = (dcifimemload_19 & ((\Mux51~16_combout  & ((\Mux51~18_combout ))) # (!\Mux51~16_combout  & (\Mux51~11_combout )))) # (!dcifimemload_19 & (((\Mux51~16_combout ))))

	.dataa(\Mux51~11_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux51~18_combout ),
	.datad(\Mux51~16_combout ),
	.cin(gnd),
	.combout(Mux511),
	.cout());
// synopsys translate_off
defparam \Mux51~19 .lut_mask = 16'hF388;
defparam \Mux51~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N30
cycloneive_lcell_comb \Mux19~20 (
// Equation(s):
// Mux19 = (dcifimemload_25 & (\Mux19~9_combout )) # (!dcifimemload_25 & ((\Mux19~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux19~9_combout ),
	.datad(\Mux19~19_combout ),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~20 .lut_mask = 16'hF3C0;
defparam \Mux19~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N12
cycloneive_lcell_comb \Mux52~9 (
// Equation(s):
// Mux52 = (dcifimemload_16 & ((\Mux52~6_combout  & (\Mux52~8_combout )) # (!\Mux52~6_combout  & ((\Mux52~1_combout ))))) # (!dcifimemload_16 & (((\Mux52~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux52~8_combout ),
	.datac(\Mux52~1_combout ),
	.datad(\Mux52~6_combout ),
	.cin(gnd),
	.combout(Mux52),
	.cout());
// synopsys translate_off
defparam \Mux52~9 .lut_mask = 16'hDDA0;
defparam \Mux52~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N8
cycloneive_lcell_comb \Mux52~19 (
// Equation(s):
// Mux521 = (dcifimemload_18 & ((\Mux52~16_combout  & (\Mux52~18_combout )) # (!\Mux52~16_combout  & ((\Mux52~11_combout ))))) # (!dcifimemload_18 & (((\Mux52~16_combout ))))

	.dataa(\Mux52~18_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux52~16_combout ),
	.datad(\Mux52~11_combout ),
	.cin(gnd),
	.combout(Mux521),
	.cout());
// synopsys translate_off
defparam \Mux52~19 .lut_mask = 16'hBCB0;
defparam \Mux52~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N18
cycloneive_lcell_comb \Mux20~20 (
// Equation(s):
// Mux20 = (dcifimemload_25 & ((\Mux20~9_combout ))) # (!dcifimemload_25 & (\Mux20~19_combout ))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux20~19_combout ),
	.datad(\Mux20~9_combout ),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~20 .lut_mask = 16'hFC30;
defparam \Mux20~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N10
cycloneive_lcell_comb \Mux53~9 (
// Equation(s):
// Mux53 = (dcifimemload_16 & ((\Mux53~6_combout  & (\Mux53~8_combout )) # (!\Mux53~6_combout  & ((\Mux53~1_combout ))))) # (!dcifimemload_16 & (((\Mux53~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux53~8_combout ),
	.datac(\Mux53~6_combout ),
	.datad(\Mux53~1_combout ),
	.cin(gnd),
	.combout(Mux53),
	.cout());
// synopsys translate_off
defparam \Mux53~9 .lut_mask = 16'hDAD0;
defparam \Mux53~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N30
cycloneive_lcell_comb \Mux53~19 (
// Equation(s):
// Mux531 = (dcifimemload_19 & ((\Mux53~16_combout  & (\Mux53~18_combout )) # (!\Mux53~16_combout  & ((\Mux53~11_combout ))))) # (!dcifimemload_19 & (((\Mux53~16_combout ))))

	.dataa(\Mux53~18_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux53~11_combout ),
	.datad(\Mux53~16_combout ),
	.cin(gnd),
	.combout(Mux531),
	.cout());
// synopsys translate_off
defparam \Mux53~19 .lut_mask = 16'hBBC0;
defparam \Mux53~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N22
cycloneive_lcell_comb \Mux21~20 (
// Equation(s):
// Mux21 = (dcifimemload_25 & (\Mux21~9_combout )) # (!dcifimemload_25 & ((\Mux21~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux21~9_combout ),
	.datad(\Mux21~19_combout ),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~20 .lut_mask = 16'hF3C0;
defparam \Mux21~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N6
cycloneive_lcell_comb \Mux54~9 (
// Equation(s):
// Mux54 = (dcifimemload_16 & ((\Mux54~6_combout  & ((\Mux54~8_combout ))) # (!\Mux54~6_combout  & (\Mux54~1_combout )))) # (!dcifimemload_16 & (((\Mux54~6_combout ))))

	.dataa(\Mux54~1_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux54~6_combout ),
	.datad(\Mux54~8_combout ),
	.cin(gnd),
	.combout(Mux54),
	.cout());
// synopsys translate_off
defparam \Mux54~9 .lut_mask = 16'hF838;
defparam \Mux54~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N14
cycloneive_lcell_comb \Mux54~19 (
// Equation(s):
// Mux541 = (dcifimemload_18 & ((\Mux54~16_combout  & (\Mux54~18_combout )) # (!\Mux54~16_combout  & ((\Mux54~11_combout ))))) # (!dcifimemload_18 & (((\Mux54~16_combout ))))

	.dataa(\Mux54~18_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux54~11_combout ),
	.datad(\Mux54~16_combout ),
	.cin(gnd),
	.combout(Mux541),
	.cout());
// synopsys translate_off
defparam \Mux54~19 .lut_mask = 16'hBBC0;
defparam \Mux54~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N6
cycloneive_lcell_comb \Mux22~20 (
// Equation(s):
// Mux22 = (dcifimemload_25 & (\Mux22~9_combout )) # (!dcifimemload_25 & ((\Mux22~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux22~9_combout ),
	.datad(\Mux22~19_combout ),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~20 .lut_mask = 16'hF5A0;
defparam \Mux22~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N26
cycloneive_lcell_comb \Mux55~9 (
// Equation(s):
// Mux55 = (dcifimemload_16 & ((\Mux55~6_combout  & ((\Mux55~8_combout ))) # (!\Mux55~6_combout  & (\Mux55~1_combout )))) # (!dcifimemload_16 & (\Mux55~6_combout ))

	.dataa(dcifimemload_16),
	.datab(\Mux55~6_combout ),
	.datac(\Mux55~1_combout ),
	.datad(\Mux55~8_combout ),
	.cin(gnd),
	.combout(Mux55),
	.cout());
// synopsys translate_off
defparam \Mux55~9 .lut_mask = 16'hEC64;
defparam \Mux55~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N16
cycloneive_lcell_comb \Mux55~19 (
// Equation(s):
// Mux551 = (dcifimemload_19 & ((\Mux55~16_combout  & ((\Mux55~18_combout ))) # (!\Mux55~16_combout  & (\Mux55~11_combout )))) # (!dcifimemload_19 & (((\Mux55~16_combout ))))

	.dataa(\Mux55~11_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux55~18_combout ),
	.datad(\Mux55~16_combout ),
	.cin(gnd),
	.combout(Mux551),
	.cout());
// synopsys translate_off
defparam \Mux55~19 .lut_mask = 16'hF388;
defparam \Mux55~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N14
cycloneive_lcell_comb \Mux23~20 (
// Equation(s):
// Mux23 = (dcifimemload_25 & (\Mux23~9_combout )) # (!dcifimemload_25 & ((\Mux23~19_combout )))

	.dataa(dcifimemload_25),
	.datab(\Mux23~9_combout ),
	.datac(gnd),
	.datad(\Mux23~19_combout ),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~20 .lut_mask = 16'hDD88;
defparam \Mux23~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N10
cycloneive_lcell_comb \Mux56~9 (
// Equation(s):
// Mux56 = (dcifimemload_16 & ((\Mux56~6_combout  & ((\Mux56~8_combout ))) # (!\Mux56~6_combout  & (\Mux56~1_combout )))) # (!dcifimemload_16 & (((\Mux56~6_combout ))))

	.dataa(\Mux56~1_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux56~6_combout ),
	.datad(\Mux56~8_combout ),
	.cin(gnd),
	.combout(Mux56),
	.cout());
// synopsys translate_off
defparam \Mux56~9 .lut_mask = 16'hF838;
defparam \Mux56~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N2
cycloneive_lcell_comb \Mux56~19 (
// Equation(s):
// Mux561 = (dcifimemload_18 & ((\Mux56~16_combout  & (\Mux56~18_combout )) # (!\Mux56~16_combout  & ((\Mux56~11_combout ))))) # (!dcifimemload_18 & (((\Mux56~16_combout ))))

	.dataa(\Mux56~18_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux56~11_combout ),
	.datad(\Mux56~16_combout ),
	.cin(gnd),
	.combout(Mux561),
	.cout());
// synopsys translate_off
defparam \Mux56~19 .lut_mask = 16'hBBC0;
defparam \Mux56~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N26
cycloneive_lcell_comb \Mux24~20 (
// Equation(s):
// Mux24 = (dcifimemload_25 & ((\Mux24~9_combout ))) # (!dcifimemload_25 & (\Mux24~19_combout ))

	.dataa(gnd),
	.datab(\Mux24~19_combout ),
	.datac(dcifimemload_25),
	.datad(\Mux24~9_combout ),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~20 .lut_mask = 16'hFC0C;
defparam \Mux24~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N2
cycloneive_lcell_comb \Mux57~9 (
// Equation(s):
// Mux57 = (dcifimemload_16 & ((\Mux57~6_combout  & ((\Mux57~8_combout ))) # (!\Mux57~6_combout  & (\Mux57~1_combout )))) # (!dcifimemload_16 & (((\Mux57~6_combout ))))

	.dataa(\Mux57~1_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux57~8_combout ),
	.datad(\Mux57~6_combout ),
	.cin(gnd),
	.combout(Mux57),
	.cout());
// synopsys translate_off
defparam \Mux57~9 .lut_mask = 16'hF388;
defparam \Mux57~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N26
cycloneive_lcell_comb \Mux57~19 (
// Equation(s):
// Mux571 = (dcifimemload_19 & ((\Mux57~16_combout  & (\Mux57~18_combout )) # (!\Mux57~16_combout  & ((\Mux57~11_combout ))))) # (!dcifimemload_19 & (((\Mux57~16_combout ))))

	.dataa(\Mux57~18_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux57~11_combout ),
	.datad(\Mux57~16_combout ),
	.cin(gnd),
	.combout(Mux571),
	.cout());
// synopsys translate_off
defparam \Mux57~19 .lut_mask = 16'hBBC0;
defparam \Mux57~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N14
cycloneive_lcell_comb \Mux25~20 (
// Equation(s):
// Mux25 = (dcifimemload_25 & (\Mux25~9_combout )) # (!dcifimemload_25 & ((\Mux25~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux25~9_combout ),
	.datad(\Mux25~19_combout ),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~20 .lut_mask = 16'hF5A0;
defparam \Mux25~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N30
cycloneive_lcell_comb \Mux58~9 (
// Equation(s):
// Mux58 = (dcifimemload_16 & ((\Mux58~6_combout  & (\Mux58~8_combout )) # (!\Mux58~6_combout  & ((\Mux58~1_combout ))))) # (!dcifimemload_16 & (((\Mux58~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux58~8_combout ),
	.datac(\Mux58~1_combout ),
	.datad(\Mux58~6_combout ),
	.cin(gnd),
	.combout(Mux58),
	.cout());
// synopsys translate_off
defparam \Mux58~9 .lut_mask = 16'hDDA0;
defparam \Mux58~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N18
cycloneive_lcell_comb \Mux58~19 (
// Equation(s):
// Mux581 = (dcifimemload_18 & ((\Mux58~16_combout  & (\Mux58~18_combout )) # (!\Mux58~16_combout  & ((\Mux58~11_combout ))))) # (!dcifimemload_18 & (((\Mux58~16_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux58~18_combout ),
	.datac(\Mux58~16_combout ),
	.datad(\Mux58~11_combout ),
	.cin(gnd),
	.combout(Mux581),
	.cout());
// synopsys translate_off
defparam \Mux58~19 .lut_mask = 16'hDAD0;
defparam \Mux58~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N12
cycloneive_lcell_comb \Mux26~20 (
// Equation(s):
// Mux26 = (dcifimemload_25 & ((\Mux26~9_combout ))) # (!dcifimemload_25 & (\Mux26~19_combout ))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux26~19_combout ),
	.datad(\Mux26~9_combout ),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~20 .lut_mask = 16'hFC30;
defparam \Mux26~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N30
cycloneive_lcell_comb \Mux59~9 (
// Equation(s):
// Mux59 = (dcifimemload_16 & ((\Mux59~6_combout  & (\Mux59~8_combout )) # (!\Mux59~6_combout  & ((\Mux59~1_combout ))))) # (!dcifimemload_16 & (((\Mux59~6_combout ))))

	.dataa(\Mux59~8_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux59~6_combout ),
	.datad(\Mux59~1_combout ),
	.cin(gnd),
	.combout(Mux59),
	.cout());
// synopsys translate_off
defparam \Mux59~9 .lut_mask = 16'hBCB0;
defparam \Mux59~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N18
cycloneive_lcell_comb \Mux59~19 (
// Equation(s):
// Mux591 = (dcifimemload_19 & ((\Mux59~16_combout  & (\Mux59~18_combout )) # (!\Mux59~16_combout  & ((\Mux59~11_combout ))))) # (!dcifimemload_19 & (((\Mux59~16_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux59~18_combout ),
	.datac(\Mux59~11_combout ),
	.datad(\Mux59~16_combout ),
	.cin(gnd),
	.combout(Mux591),
	.cout());
// synopsys translate_off
defparam \Mux59~19 .lut_mask = 16'hDDA0;
defparam \Mux59~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N0
cycloneive_lcell_comb \Mux27~20 (
// Equation(s):
// Mux27 = (dcifimemload_25 & (\Mux27~9_combout )) # (!dcifimemload_25 & ((\Mux27~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux27~9_combout ),
	.datad(\Mux27~19_combout ),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~20 .lut_mask = 16'hF5A0;
defparam \Mux27~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N10
cycloneive_lcell_comb \Mux60~9 (
// Equation(s):
// Mux60 = (dcifimemload_16 & ((\Mux60~6_combout  & ((\Mux60~8_combout ))) # (!\Mux60~6_combout  & (\Mux60~1_combout )))) # (!dcifimemload_16 & (((\Mux60~6_combout ))))

	.dataa(\Mux60~1_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux60~6_combout ),
	.datad(\Mux60~8_combout ),
	.cin(gnd),
	.combout(Mux60),
	.cout());
// synopsys translate_off
defparam \Mux60~9 .lut_mask = 16'hF838;
defparam \Mux60~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N2
cycloneive_lcell_comb \Mux60~19 (
// Equation(s):
// Mux601 = (dcifimemload_18 & ((\Mux60~16_combout  & (\Mux60~18_combout )) # (!\Mux60~16_combout  & ((\Mux60~11_combout ))))) # (!dcifimemload_18 & (((\Mux60~16_combout ))))

	.dataa(\Mux60~18_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux60~11_combout ),
	.datad(\Mux60~16_combout ),
	.cin(gnd),
	.combout(Mux601),
	.cout());
// synopsys translate_off
defparam \Mux60~19 .lut_mask = 16'hBBC0;
defparam \Mux60~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N0
cycloneive_lcell_comb \Mux28~20 (
// Equation(s):
// Mux28 = (dcifimemload_25 & (\Mux28~9_combout )) # (!dcifimemload_25 & ((\Mux28~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux28~9_combout ),
	.datad(\Mux28~19_combout ),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~20 .lut_mask = 16'hF3C0;
defparam \Mux28~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N8
cycloneive_lcell_comb \Mux61~9 (
// Equation(s):
// Mux61 = (dcifimemload_16 & ((\Mux61~6_combout  & (\Mux61~8_combout )) # (!\Mux61~6_combout  & ((\Mux61~1_combout ))))) # (!dcifimemload_16 & (\Mux61~6_combout ))

	.dataa(dcifimemload_16),
	.datab(\Mux61~6_combout ),
	.datac(\Mux61~8_combout ),
	.datad(\Mux61~1_combout ),
	.cin(gnd),
	.combout(Mux61),
	.cout());
// synopsys translate_off
defparam \Mux61~9 .lut_mask = 16'hE6C4;
defparam \Mux61~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N20
cycloneive_lcell_comb \Mux61~19 (
// Equation(s):
// Mux611 = (dcifimemload_19 & ((\Mux61~16_combout  & (\Mux61~18_combout )) # (!\Mux61~16_combout  & ((\Mux61~11_combout ))))) # (!dcifimemload_19 & (((\Mux61~16_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux61~18_combout ),
	.datac(\Mux61~16_combout ),
	.datad(\Mux61~11_combout ),
	.cin(gnd),
	.combout(Mux611),
	.cout());
// synopsys translate_off
defparam \Mux61~19 .lut_mask = 16'hDAD0;
defparam \Mux61~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N22
cycloneive_lcell_comb \Mux29~20 (
// Equation(s):
// Mux29 = (dcifimemload_25 & (\Mux29~9_combout )) # (!dcifimemload_25 & ((\Mux29~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux29~9_combout ),
	.datad(\Mux29~19_combout ),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~20 .lut_mask = 16'hF3C0;
defparam \Mux29~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N26
cycloneive_lcell_comb \Mux62~9 (
// Equation(s):
// Mux62 = (dcifimemload_16 & ((\Mux62~6_combout  & ((\Mux62~8_combout ))) # (!\Mux62~6_combout  & (\Mux62~1_combout )))) # (!dcifimemload_16 & (\Mux62~6_combout ))

	.dataa(dcifimemload_16),
	.datab(\Mux62~6_combout ),
	.datac(\Mux62~1_combout ),
	.datad(\Mux62~8_combout ),
	.cin(gnd),
	.combout(Mux62),
	.cout());
// synopsys translate_off
defparam \Mux62~9 .lut_mask = 16'hEC64;
defparam \Mux62~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N0
cycloneive_lcell_comb \Mux62~19 (
// Equation(s):
// Mux621 = (dcifimemload_18 & ((\Mux62~16_combout  & ((\Mux62~18_combout ))) # (!\Mux62~16_combout  & (\Mux62~11_combout )))) # (!dcifimemload_18 & (((\Mux62~16_combout ))))

	.dataa(\Mux62~11_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux62~18_combout ),
	.datad(\Mux62~16_combout ),
	.cin(gnd),
	.combout(Mux621),
	.cout());
// synopsys translate_off
defparam \Mux62~19 .lut_mask = 16'hF388;
defparam \Mux62~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N14
cycloneive_lcell_comb \Mux31~20 (
// Equation(s):
// Mux31 = (dcifimemload_25 & (\Mux31~9_combout )) # (!dcifimemload_25 & ((\Mux31~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux31~9_combout ),
	.datad(\Mux31~19_combout ),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux31~20 .lut_mask = 16'hF3C0;
defparam \Mux31~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N8
cycloneive_lcell_comb \Mux32~9 (
// Equation(s):
// Mux32 = (dcifimemload_18 & ((\Mux32~6_combout  & (\Mux32~8_combout )) # (!\Mux32~6_combout  & ((\Mux32~1_combout ))))) # (!dcifimemload_18 & (((\Mux32~6_combout ))))

	.dataa(\Mux32~8_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux32~1_combout ),
	.datad(\Mux32~6_combout ),
	.cin(gnd),
	.combout(Mux32),
	.cout());
// synopsys translate_off
defparam \Mux32~9 .lut_mask = 16'hBBC0;
defparam \Mux32~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N14
cycloneive_lcell_comb \Mux32~19 (
// Equation(s):
// Mux321 = (dcifimemload_16 & ((\Mux32~16_combout  & (\Mux32~18_combout )) # (!\Mux32~16_combout  & ((\Mux32~11_combout ))))) # (!dcifimemload_16 & (((\Mux32~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux32~18_combout ),
	.datac(\Mux32~11_combout ),
	.datad(\Mux32~16_combout ),
	.cin(gnd),
	.combout(Mux321),
	.cout());
// synopsys translate_off
defparam \Mux32~19 .lut_mask = 16'hDDA0;
defparam \Mux32~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N0
cycloneive_lcell_comb \Mux0~20 (
// Equation(s):
// Mux0 = (dcifimemload_25 & ((\Mux0~9_combout ))) # (!dcifimemload_25 & (\Mux0~19_combout ))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux0~19_combout ),
	.datad(\Mux0~9_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~20 .lut_mask = 16'hFC30;
defparam \Mux0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N16
cycloneive_lcell_comb \regs~4 (
// Equation(s):
// \regs~4_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_01)) # (!cuifRegSel_0 & ((Mux312)))))

	.dataa(cuifRegSel_0),
	.datab(cuifRegSel_11),
	.datac(ramiframload_0),
	.datad(Mux311),
	.cin(gnd),
	.combout(\regs~4_combout ),
	.cout());
// synopsys translate_off
defparam \regs~4 .lut_mask = 16'h3120;
defparam \regs~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N22
cycloneive_lcell_comb \regs~64 (
// Equation(s):
// \regs~64_combout  = (!dcifimemload_31 & (!dcifimemload_30 & (cuifRegSel_1 & !cuifRegSel_0)))

	.dataa(dcifimemload_31),
	.datab(dcifimemload_30),
	.datac(cuifRegSel_1),
	.datad(cuifRegSel_0),
	.cin(gnd),
	.combout(\regs~64_combout ),
	.cout());
// synopsys translate_off
defparam \regs~64 .lut_mask = 16'h0010;
defparam \regs~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N20
cycloneive_lcell_comb \regs~5 (
// Equation(s):
// \regs~5_combout  = (!\Equal0~1_combout  & ((\regs~4_combout ) # ((PC_0 & \regs~64_combout ))))

	.dataa(\Equal0~1_combout ),
	.datab(\regs~4_combout ),
	.datac(PC_0),
	.datad(\regs~64_combout ),
	.cin(gnd),
	.combout(\regs~5_combout ),
	.cout());
// synopsys translate_off
defparam \regs~5 .lut_mask = 16'h5444;
defparam \regs~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N20
cycloneive_lcell_comb \regs[20][0]~feeder (
// Equation(s):
// \regs[20][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~5_combout ),
	.cin(gnd),
	.combout(\regs[20][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][0]~feeder .lut_mask = 16'hFF00;
defparam \regs[20][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N18
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!\Selector67~0_combout  & !\Selector68~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector67),
	.datad(Selector68),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h000F;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N22
cycloneive_lcell_comb \Decoder0~12 (
// Equation(s):
// \Decoder0~12_combout  = (!dcifimemload_30 & (\Equal0~0_combout  & ((Selector4) # (Selector41))))

	.dataa(dcifimemload_30),
	.datab(Selector4),
	.datac(\Equal0~0_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Decoder0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~12 .lut_mask = 16'h5040;
defparam \Decoder0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N26
cycloneive_lcell_comb \Decoder0~13 (
// Equation(s):
// \Decoder0~13_combout  = (\Selector64~0_combout  & (!\Selector65~0_combout  & (\Selector66~0_combout  & \Decoder0~12_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~13 .lut_mask = 16'h2000;
defparam \Decoder0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N21
dffeas \regs[20][0] (
	.clk(CLK),
	.d(\regs[20][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][0] .is_wysiwyg = "true";
defparam \regs[20][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N8
cycloneive_lcell_comb \Decoder0~16 (
// Equation(s):
// \Decoder0~16_combout  = (\Decoder0~12_combout  & (\Selector65~0_combout  & (\Selector64~0_combout  & \Selector66~0_combout )))

	.dataa(\Decoder0~12_combout ),
	.datab(Selector65),
	.datac(Selector64),
	.datad(Selector66),
	.cin(gnd),
	.combout(\Decoder0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~16 .lut_mask = 16'h8000;
defparam \Decoder0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N27
dffeas \regs[28][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][0] .is_wysiwyg = "true";
defparam \regs[28][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N16
cycloneive_lcell_comb \regs[24][0]~feeder (
// Equation(s):
// \regs[24][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[24][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][0]~feeder .lut_mask = 16'hF0F0;
defparam \regs[24][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N20
cycloneive_lcell_comb \Decoder0~14 (
// Equation(s):
// \Decoder0~14_combout  = (\Decoder0~12_combout  & (\Selector65~0_combout  & (\Selector64~0_combout  & !\Selector66~0_combout )))

	.dataa(\Decoder0~12_combout ),
	.datab(Selector65),
	.datac(Selector64),
	.datad(Selector66),
	.cin(gnd),
	.combout(\Decoder0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~14 .lut_mask = 16'h0080;
defparam \Decoder0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N17
dffeas \regs[24][0] (
	.clk(CLK),
	.d(\regs[24][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][0] .is_wysiwyg = "true";
defparam \regs[24][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N26
cycloneive_lcell_comb \Decoder0~15 (
// Equation(s):
// \Decoder0~15_combout  = (\Decoder0~12_combout  & (!\Selector65~0_combout  & (\Selector64~0_combout  & !\Selector66~0_combout )))

	.dataa(\Decoder0~12_combout ),
	.datab(Selector65),
	.datac(Selector64),
	.datad(Selector66),
	.cin(gnd),
	.combout(\Decoder0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~15 .lut_mask = 16'h0020;
defparam \Decoder0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N21
dffeas \regs[16][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][0] .is_wysiwyg = "true";
defparam \regs[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N20
cycloneive_lcell_comb \Mux63~4 (
// Equation(s):
// \Mux63~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[24][0]~q )) # (!dcifimemload_19 & ((\regs[16][0]~q )))))

	.dataa(dcifimemload_18),
	.datab(\regs[24][0]~q ),
	.datac(\regs[16][0]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux63~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~4 .lut_mask = 16'hEE50;
defparam \Mux63~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N26
cycloneive_lcell_comb \Mux63~5 (
// Equation(s):
// \Mux63~5_combout  = (dcifimemload_18 & ((\Mux63~4_combout  & ((\regs[28][0]~q ))) # (!\Mux63~4_combout  & (\regs[20][0]~q )))) # (!dcifimemload_18 & (((\Mux63~4_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[20][0]~q ),
	.datac(\regs[28][0]~q ),
	.datad(\Mux63~4_combout ),
	.cin(gnd),
	.combout(\Mux63~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~5 .lut_mask = 16'hF588;
defparam \Mux63~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N26
cycloneive_lcell_comb \Decoder0~7 (
// Equation(s):
// \Decoder0~7_combout  = (\Selector67~0_combout  & (!\Selector68~1_combout  & Selector42))

	.dataa(Selector67),
	.datab(gnd),
	.datac(Selector68),
	.datad(Selector42),
	.cin(gnd),
	.combout(\Decoder0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~7 .lut_mask = 16'h0A00;
defparam \Decoder0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N30
cycloneive_lcell_comb \Decoder0~10 (
// Equation(s):
// \Decoder0~10_combout  = (\Selector64~0_combout  & (!\Selector65~0_combout  & (!\Selector66~0_combout  & \Decoder0~7_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\Decoder0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~10 .lut_mask = 16'h0200;
defparam \Decoder0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N5
dffeas \regs[18][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][0] .is_wysiwyg = "true";
defparam \regs[18][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N4
cycloneive_lcell_comb \Mux63~2 (
// Equation(s):
// \Mux63~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[26][0]~q )) # (!dcifimemload_19 & ((\regs[18][0]~q )))))

	.dataa(\regs[26][0]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][0]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux63~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~2 .lut_mask = 16'hEE30;
defparam \Mux63~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N18
cycloneive_lcell_comb \Decoder0~11 (
// Equation(s):
// \Decoder0~11_combout  = (\Selector64~0_combout  & (\Selector66~0_combout  & (\Selector65~0_combout  & \Decoder0~7_combout )))

	.dataa(Selector64),
	.datab(Selector66),
	.datac(Selector65),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\Decoder0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~11 .lut_mask = 16'h8000;
defparam \Decoder0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N15
dffeas \regs[30][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][0] .is_wysiwyg = "true";
defparam \regs[30][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N14
cycloneive_lcell_comb \Mux63~3 (
// Equation(s):
// \Mux63~3_combout  = (\Mux63~2_combout  & (((\regs[30][0]~q ) # (!dcifimemload_18)))) # (!\Mux63~2_combout  & (\regs[22][0]~q  & ((dcifimemload_18))))

	.dataa(\regs[22][0]~q ),
	.datab(\Mux63~2_combout ),
	.datac(\regs[30][0]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux63~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~3 .lut_mask = 16'hE2CC;
defparam \Mux63~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N8
cycloneive_lcell_comb \Mux63~6 (
// Equation(s):
// \Mux63~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux63~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux63~5_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux63~5_combout ),
	.datad(\Mux63~3_combout ),
	.cin(gnd),
	.combout(\Mux63~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~6 .lut_mask = 16'hBA98;
defparam \Mux63~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N10
cycloneive_lcell_comb \Decoder0~0 (
// Equation(s):
// \Decoder0~0_combout  = (\Selector68~1_combout  & (!dcifimemload_30 & ((Selector4) # (Selector41))))

	.dataa(Selector68),
	.datab(Selector4),
	.datac(dcifimemload_30),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~0 .lut_mask = 16'h0A08;
defparam \Decoder0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N0
cycloneive_lcell_comb \Decoder0~1 (
// Equation(s):
// \Decoder0~1_combout  = (\Decoder0~0_combout  & !\Selector67~0_combout )

	.dataa(gnd),
	.datab(\Decoder0~0_combout ),
	.datac(gnd),
	.datad(Selector67),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~1 .lut_mask = 16'h00CC;
defparam \Decoder0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N18
cycloneive_lcell_comb \Decoder0~2 (
// Equation(s):
// \Decoder0~2_combout  = (\Selector64~0_combout  & (\Selector65~0_combout  & (!\Selector66~0_combout  & \Decoder0~1_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~1_combout ),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~2 .lut_mask = 16'h0800;
defparam \Decoder0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N17
dffeas \regs[25][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][0] .is_wysiwyg = "true";
defparam \regs[25][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N2
cycloneive_lcell_comb \Decoder0~3 (
// Equation(s):
// \Decoder0~3_combout  = (!\Selector67~0_combout  & (\Selector66~0_combout  & \Decoder0~0_combout ))

	.dataa(Selector67),
	.datab(Selector66),
	.datac(gnd),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~3 .lut_mask = 16'h4400;
defparam \Decoder0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N12
cycloneive_lcell_comb \Decoder0~6 (
// Equation(s):
// \Decoder0~6_combout  = (\Selector65~0_combout  & (\Selector64~0_combout  & \Decoder0~3_combout ))

	.dataa(Selector65),
	.datab(Selector64),
	.datac(gnd),
	.datad(\Decoder0~3_combout ),
	.cin(gnd),
	.combout(\Decoder0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~6 .lut_mask = 16'h8800;
defparam \Decoder0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N19
dffeas \regs[29][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][0] .is_wysiwyg = "true";
defparam \regs[29][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N16
cycloneive_lcell_comb \regs[17][0]~feeder (
// Equation(s):
// \regs[17][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~5_combout ),
	.cin(gnd),
	.combout(\regs[17][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][0]~feeder .lut_mask = 16'hFF00;
defparam \regs[17][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N24
cycloneive_lcell_comb \Decoder0~5 (
// Equation(s):
// \Decoder0~5_combout  = (\Selector64~0_combout  & (!\Selector65~0_combout  & (!\Selector66~0_combout  & \Decoder0~1_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~1_combout ),
	.cin(gnd),
	.combout(\Decoder0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~5 .lut_mask = 16'h0200;
defparam \Decoder0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N17
dffeas \regs[17][0] (
	.clk(CLK),
	.d(\regs[17][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][0] .is_wysiwyg = "true";
defparam \regs[17][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N24
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (dcifimemload_18 & ((\regs[21][0]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[17][0]~q  & !dcifimemload_19))))

	.dataa(\regs[21][0]~q ),
	.datab(\regs[17][0]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hF0AC;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N18
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (dcifimemload_19 & ((\Mux63~0_combout  & ((\regs[29][0]~q ))) # (!\Mux63~0_combout  & (\regs[25][0]~q )))) # (!dcifimemload_19 & (((\Mux63~0_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[25][0]~q ),
	.datac(\regs[29][0]~q ),
	.datad(\Mux63~0_combout ),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hF588;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N0
cycloneive_lcell_comb \Decoder0~17 (
// Equation(s):
// \Decoder0~17_combout  = (\Selector67~0_combout  & \Decoder0~0_combout )

	.dataa(Selector67),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~17 .lut_mask = 16'hAA00;
defparam \Decoder0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N16
cycloneive_lcell_comb \Decoder0~18 (
// Equation(s):
// \Decoder0~18_combout  = (\Selector65~0_combout  & (\Selector64~0_combout  & (\Decoder0~17_combout  & !\Selector66~0_combout )))

	.dataa(Selector65),
	.datab(Selector64),
	.datac(\Decoder0~17_combout ),
	.datad(Selector66),
	.cin(gnd),
	.combout(\Decoder0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~18 .lut_mask = 16'h0080;
defparam \Decoder0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N9
dffeas \regs[27][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][0] .is_wysiwyg = "true";
defparam \regs[27][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N8
cycloneive_lcell_comb \regs[31][0]~feeder (
// Equation(s):
// \regs[31][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[31][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][0]~feeder .lut_mask = 16'hF0F0;
defparam \regs[31][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N22
cycloneive_lcell_comb \Decoder0~21 (
// Equation(s):
// \Decoder0~21_combout  = (\Selector65~0_combout  & (\Selector64~0_combout  & (\Decoder0~17_combout  & \Selector66~0_combout )))

	.dataa(Selector65),
	.datab(Selector64),
	.datac(\Decoder0~17_combout ),
	.datad(Selector66),
	.cin(gnd),
	.combout(\Decoder0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~21 .lut_mask = 16'h8000;
defparam \Decoder0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N9
dffeas \regs[31][0] (
	.clk(CLK),
	.d(\regs[31][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][0] .is_wysiwyg = "true";
defparam \regs[31][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N4
cycloneive_lcell_comb \regs[23][0]~feeder (
// Equation(s):
// \regs[23][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[23][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][0]~feeder .lut_mask = 16'hF0F0;
defparam \regs[23][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N18
cycloneive_lcell_comb \Decoder0~19 (
// Equation(s):
// \Decoder0~19_combout  = (!\Selector65~0_combout  & (\Selector64~0_combout  & (\Decoder0~17_combout  & \Selector66~0_combout )))

	.dataa(Selector65),
	.datab(Selector64),
	.datac(\Decoder0~17_combout ),
	.datad(Selector66),
	.cin(gnd),
	.combout(\Decoder0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~19 .lut_mask = 16'h4000;
defparam \Decoder0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N5
dffeas \regs[23][0] (
	.clk(CLK),
	.d(\regs[23][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][0] .is_wysiwyg = "true";
defparam \regs[23][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N2
cycloneive_lcell_comb \Mux63~7 (
// Equation(s):
// \Mux63~7_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\regs[23][0]~q ))) # (!dcifimemload_18 & (\regs[19][0]~q ))))

	.dataa(\regs[19][0]~q ),
	.datab(\regs[23][0]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux63~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~7 .lut_mask = 16'hFC0A;
defparam \Mux63~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N14
cycloneive_lcell_comb \Mux63~8 (
// Equation(s):
// \Mux63~8_combout  = (dcifimemload_19 & ((\Mux63~7_combout  & ((\regs[31][0]~q ))) # (!\Mux63~7_combout  & (\regs[27][0]~q )))) # (!dcifimemload_19 & (((\Mux63~7_combout ))))

	.dataa(\regs[27][0]~q ),
	.datab(\regs[31][0]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux63~7_combout ),
	.cin(gnd),
	.combout(\Mux63~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~8 .lut_mask = 16'hCFA0;
defparam \Mux63~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N30
cycloneive_lcell_comb \regs[9][0]~feeder (
// Equation(s):
// \regs[9][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~5_combout ),
	.cin(gnd),
	.combout(\regs[9][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][0]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N12
cycloneive_lcell_comb \Decoder0~22 (
// Equation(s):
// \Decoder0~22_combout  = (!\Selector64~0_combout  & (!\Selector66~0_combout  & (\Selector65~0_combout  & \Decoder0~1_combout )))

	.dataa(Selector64),
	.datab(Selector66),
	.datac(Selector65),
	.datad(\Decoder0~1_combout ),
	.cin(gnd),
	.combout(\Decoder0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~22 .lut_mask = 16'h1000;
defparam \Decoder0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N31
dffeas \regs[9][0] (
	.clk(CLK),
	.d(\regs[9][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][0] .is_wysiwyg = "true";
defparam \regs[9][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N12
cycloneive_lcell_comb \Decoder0~25 (
// Equation(s):
// \Decoder0~25_combout  = (!\Selector64~0_combout  & (\Decoder0~0_combout  & \Selector67~0_combout ))

	.dataa(Selector64),
	.datab(\Decoder0~0_combout ),
	.datac(Selector67),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~25 .lut_mask = 16'h4040;
defparam \Decoder0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N8
cycloneive_lcell_comb \Decoder0~26 (
// Equation(s):
// \Decoder0~26_combout  = (!\Selector66~0_combout  & (\Selector65~0_combout  & \Decoder0~25_combout ))

	.dataa(Selector66),
	.datab(Selector65),
	.datac(gnd),
	.datad(\Decoder0~25_combout ),
	.cin(gnd),
	.combout(\Decoder0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~26 .lut_mask = 16'h4400;
defparam \Decoder0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N7
dffeas \regs[11][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][0] .is_wysiwyg = "true";
defparam \regs[11][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N28
cycloneive_lcell_comb \Decoder0~24 (
// Equation(s):
// \Decoder0~24_combout  = (!\Selector64~0_combout  & (\Selector65~0_combout  & (!\Selector66~0_combout  & \Decoder0~12_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~24 .lut_mask = 16'h0400;
defparam \Decoder0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N25
dffeas \regs[8][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][0] .is_wysiwyg = "true";
defparam \regs[8][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N0
cycloneive_lcell_comb \Decoder0~23 (
// Equation(s):
// \Decoder0~23_combout  = (!\Selector64~0_combout  & (\Selector65~0_combout  & (!\Selector66~0_combout  & \Decoder0~7_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\Decoder0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~23 .lut_mask = 16'h0400;
defparam \Decoder0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N21
dffeas \regs[10][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][0] .is_wysiwyg = "true";
defparam \regs[10][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N24
cycloneive_lcell_comb \Mux63~10 (
// Equation(s):
// \Mux63~10_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\regs[10][0]~q )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\regs[8][0]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[8][0]~q ),
	.datad(\regs[10][0]~q ),
	.cin(gnd),
	.combout(\Mux63~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~10 .lut_mask = 16'hBA98;
defparam \Mux63~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N6
cycloneive_lcell_comb \Mux63~11 (
// Equation(s):
// \Mux63~11_combout  = (dcifimemload_16 & ((\Mux63~10_combout  & ((\regs[11][0]~q ))) # (!\Mux63~10_combout  & (\regs[9][0]~q )))) # (!dcifimemload_16 & (((\Mux63~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][0]~q ),
	.datac(\regs[11][0]~q ),
	.datad(\Mux63~10_combout ),
	.cin(gnd),
	.combout(\Mux63~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~11 .lut_mask = 16'hF588;
defparam \Mux63~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N18
cycloneive_lcell_comb \Decoder0~34 (
// Equation(s):
// \Decoder0~34_combout  = (!\Selector64~0_combout  & (\Selector65~0_combout  & (\Selector66~0_combout  & \Decoder0~7_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\Decoder0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~34 .lut_mask = 16'h4000;
defparam \Decoder0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N27
dffeas \regs[14][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][0] .is_wysiwyg = "true";
defparam \regs[14][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N4
cycloneive_lcell_comb \Decoder0~37 (
// Equation(s):
// \Decoder0~37_combout  = (\Selector66~0_combout  & (\Selector65~0_combout  & \Decoder0~25_combout ))

	.dataa(Selector66),
	.datab(Selector65),
	.datac(gnd),
	.datad(\Decoder0~25_combout ),
	.cin(gnd),
	.combout(\Decoder0~37_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~37 .lut_mask = 16'h8800;
defparam \Decoder0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y31_N3
dffeas \regs[15][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][0] .is_wysiwyg = "true";
defparam \regs[15][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N30
cycloneive_lcell_comb \Decoder0~36 (
// Equation(s):
// \Decoder0~36_combout  = (\Selector65~0_combout  & (\Decoder0~12_combout  & (\Selector66~0_combout  & !\Selector64~0_combout )))

	.dataa(Selector65),
	.datab(\Decoder0~12_combout ),
	.datac(Selector66),
	.datad(Selector64),
	.cin(gnd),
	.combout(\Decoder0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~36 .lut_mask = 16'h0080;
defparam \Decoder0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y31_N13
dffeas \regs[12][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][0] .is_wysiwyg = "true";
defparam \regs[12][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N12
cycloneive_lcell_comb \Mux63~17 (
// Equation(s):
// \Mux63~17_combout  = (dcifimemload_16 & ((\regs[13][0]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[12][0]~q  & !dcifimemload_17))))

	.dataa(\regs[13][0]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[12][0]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux63~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~17 .lut_mask = 16'hCCB8;
defparam \Mux63~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N2
cycloneive_lcell_comb \Mux63~18 (
// Equation(s):
// \Mux63~18_combout  = (dcifimemload_17 & ((\Mux63~17_combout  & ((\regs[15][0]~q ))) # (!\Mux63~17_combout  & (\regs[14][0]~q )))) # (!dcifimemload_17 & (((\Mux63~17_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[14][0]~q ),
	.datac(\regs[15][0]~q ),
	.datad(\Mux63~17_combout ),
	.cin(gnd),
	.combout(\Mux63~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~18 .lut_mask = 16'hF588;
defparam \Mux63~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \Decoder0~29 (
// Equation(s):
// \Decoder0~29_combout  = (!\Selector64~0_combout  & (!\Selector65~0_combout  & (\Selector66~0_combout  & \Decoder0~12_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~29 .lut_mask = 16'h1000;
defparam \Decoder0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N5
dffeas \regs[4][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][0] .is_wysiwyg = "true";
defparam \regs[4][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \Decoder0~28 (
// Equation(s):
// \Decoder0~28_combout  = (!\Selector64~0_combout  & (!\Selector65~0_combout  & \Decoder0~3_combout ))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(gnd),
	.datad(\Decoder0~3_combout ),
	.cin(gnd),
	.combout(\Decoder0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~28 .lut_mask = 16'h1100;
defparam \Decoder0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N19
dffeas \regs[5][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][0] .is_wysiwyg = "true";
defparam \regs[5][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N4
cycloneive_lcell_comb \Mux63~12 (
// Equation(s):
// \Mux63~12_combout  = (dcifimemload_17 & (dcifimemload_16)) # (!dcifimemload_17 & ((dcifimemload_16 & ((\regs[5][0]~q ))) # (!dcifimemload_16 & (\regs[4][0]~q ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[4][0]~q ),
	.datad(\regs[5][0]~q ),
	.cin(gnd),
	.combout(\Mux63~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~12 .lut_mask = 16'hDC98;
defparam \Mux63~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N0
cycloneive_lcell_comb \Decoder0~30 (
// Equation(s):
// \Decoder0~30_combout  = (\Selector66~0_combout  & (!\Selector65~0_combout  & \Decoder0~25_combout ))

	.dataa(Selector66),
	.datab(Selector65),
	.datac(gnd),
	.datad(\Decoder0~25_combout ),
	.cin(gnd),
	.combout(\Decoder0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~30 .lut_mask = 16'h2200;
defparam \Decoder0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N19
dffeas \regs[7][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][0] .is_wysiwyg = "true";
defparam \regs[7][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N18
cycloneive_lcell_comb \Mux63~13 (
// Equation(s):
// \Mux63~13_combout  = (\Mux63~12_combout  & (((\regs[7][0]~q ) # (!dcifimemload_17)))) # (!\Mux63~12_combout  & (\regs[6][0]~q  & ((dcifimemload_17))))

	.dataa(\regs[6][0]~q ),
	.datab(\Mux63~12_combout ),
	.datac(\regs[7][0]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux63~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~13 .lut_mask = 16'hE2CC;
defparam \Mux63~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N2
cycloneive_lcell_comb \Decoder0~31 (
// Equation(s):
// \Decoder0~31_combout  = (!\Selector64~0_combout  & (!\Selector65~0_combout  & (!\Selector66~0_combout  & \Decoder0~1_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~1_combout ),
	.cin(gnd),
	.combout(\Decoder0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~31 .lut_mask = 16'h0100;
defparam \Decoder0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N17
dffeas \regs[1][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][0] .is_wysiwyg = "true";
defparam \regs[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N24
cycloneive_lcell_comb \Decoder0~33 (
// Equation(s):
// \Decoder0~33_combout  = (!\Selector65~0_combout  & (!\Selector64~0_combout  & (\Decoder0~17_combout  & !\Selector66~0_combout )))

	.dataa(Selector65),
	.datab(Selector64),
	.datac(\Decoder0~17_combout ),
	.datad(Selector66),
	.cin(gnd),
	.combout(\Decoder0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~33 .lut_mask = 16'h0010;
defparam \Decoder0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N11
dffeas \regs[3][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][0] .is_wysiwyg = "true";
defparam \regs[3][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N10
cycloneive_lcell_comb \Mux63~14 (
// Equation(s):
// \Mux63~14_combout  = (dcifimemload_16 & ((\regs[3][0]~q ))) # (!dcifimemload_16 & (\regs[2][0]~q ))

	.dataa(\regs[2][0]~q ),
	.datab(gnd),
	.datac(\regs[3][0]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux63~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~14 .lut_mask = 16'hF0AA;
defparam \Mux63~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N16
cycloneive_lcell_comb \Mux63~15 (
// Equation(s):
// \Mux63~15_combout  = (dcifimemload_17 & (((\Mux63~14_combout )))) # (!dcifimemload_17 & (dcifimemload_16 & (\regs[1][0]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[1][0]~q ),
	.datad(\Mux63~14_combout ),
	.cin(gnd),
	.combout(\Mux63~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~15 .lut_mask = 16'hEC20;
defparam \Mux63~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N6
cycloneive_lcell_comb \Mux63~16 (
// Equation(s):
// \Mux63~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & (\Mux63~13_combout )) # (!dcifimemload_18 & ((\Mux63~15_combout )))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux63~13_combout ),
	.datad(\Mux63~15_combout ),
	.cin(gnd),
	.combout(\Mux63~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~16 .lut_mask = 16'hD9C8;
defparam \Mux63~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N20
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// \Equal0~1_combout  = (!\Selector64~0_combout  & (!\Selector66~0_combout  & (!\Selector65~0_combout  & \Equal0~0_combout )))

	.dataa(Selector64),
	.datab(Selector66),
	.datac(Selector65),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'h0100;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N6
cycloneive_lcell_comb \regs~6 (
// Equation(s):
// \regs~6_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_1)) # (!cuifRegSel_0 & ((Mux301)))))

	.dataa(cuifRegSel_0),
	.datab(ramiframload_1),
	.datac(Mux301),
	.datad(cuifRegSel_11),
	.cin(gnd),
	.combout(\regs~6_combout ),
	.cout());
// synopsys translate_off
defparam \regs~6 .lut_mask = 16'h00D8;
defparam \regs~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N6
cycloneive_lcell_comb \regs~7 (
// Equation(s):
// \regs~7_combout  = (!\Equal0~1_combout  & ((\regs~6_combout ) # ((\regs~64_combout  & PC_1))))

	.dataa(\regs~64_combout ),
	.datab(PC_1),
	.datac(\Equal0~1_combout ),
	.datad(\regs~6_combout ),
	.cin(gnd),
	.combout(\regs~7_combout ),
	.cout());
// synopsys translate_off
defparam \regs~7 .lut_mask = 16'h0F08;
defparam \regs~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N4
cycloneive_lcell_comb \regs[31][1]~feeder (
// Equation(s):
// \regs[31][1]~feeder_combout  = \regs~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[31][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][1]~feeder .lut_mask = 16'hF0F0;
defparam \regs[31][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N5
dffeas \regs[31][1] (
	.clk(CLK),
	.d(\regs[31][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][1] .is_wysiwyg = "true";
defparam \regs[31][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N10
cycloneive_lcell_comb \regs[19][1]~feeder (
// Equation(s):
// \regs[19][1]~feeder_combout  = \regs~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[19][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][1]~feeder .lut_mask = 16'hF0F0;
defparam \regs[19][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N8
cycloneive_lcell_comb \Decoder0~20 (
// Equation(s):
// \Decoder0~20_combout  = (!\Selector65~0_combout  & (\Selector64~0_combout  & (\Decoder0~17_combout  & !\Selector66~0_combout )))

	.dataa(Selector65),
	.datab(Selector64),
	.datac(\Decoder0~17_combout ),
	.datad(Selector66),
	.cin(gnd),
	.combout(\Decoder0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~20 .lut_mask = 16'h0040;
defparam \Decoder0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N11
dffeas \regs[19][1] (
	.clk(CLK),
	.d(\regs[19][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][1] .is_wysiwyg = "true";
defparam \regs[19][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N10
cycloneive_lcell_comb \Mux30~7 (
// Equation(s):
// \Mux30~7_combout  = (dcifimemload_23 & ((\regs[23][1]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[19][1]~q  & !dcifimemload_24))))

	.dataa(\regs[23][1]~q ),
	.datab(\regs[19][1]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~7 .lut_mask = 16'hF0AC;
defparam \Mux30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N8
cycloneive_lcell_comb \Mux30~8 (
// Equation(s):
// \Mux30~8_combout  = (dcifimemload_24 & ((\Mux30~7_combout  & ((\regs[31][1]~q ))) # (!\Mux30~7_combout  & (\regs[27][1]~q )))) # (!dcifimemload_24 & (((\Mux30~7_combout ))))

	.dataa(\regs[27][1]~q ),
	.datab(\regs[31][1]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux30~7_combout ),
	.cin(gnd),
	.combout(\Mux30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~8 .lut_mask = 16'hCFA0;
defparam \Mux30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N4
cycloneive_lcell_comb \regs[29][1]~feeder (
// Equation(s):
// \regs[29][1]~feeder_combout  = \regs~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[29][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][1]~feeder .lut_mask = 16'hF0F0;
defparam \regs[29][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N5
dffeas \regs[29][1] (
	.clk(CLK),
	.d(\regs[29][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][1] .is_wysiwyg = "true";
defparam \regs[29][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N26
cycloneive_lcell_comb \regs[25][1]~feeder (
// Equation(s):
// \regs[25][1]~feeder_combout  = \regs~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~7_combout ),
	.cin(gnd),
	.combout(\regs[25][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[25][1]~feeder .lut_mask = 16'hFF00;
defparam \regs[25][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N27
dffeas \regs[25][1] (
	.clk(CLK),
	.d(\regs[25][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][1] .is_wysiwyg = "true";
defparam \regs[25][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N16
cycloneive_lcell_comb \regs[21][1]~feeder (
// Equation(s):
// \regs[21][1]~feeder_combout  = \regs~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[21][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][1]~feeder .lut_mask = 16'hF0F0;
defparam \regs[21][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N26
cycloneive_lcell_comb \Decoder0~4 (
// Equation(s):
// \Decoder0~4_combout  = (!\Selector65~0_combout  & (\Selector64~0_combout  & \Decoder0~3_combout ))

	.dataa(Selector65),
	.datab(Selector64),
	.datac(gnd),
	.datad(\Decoder0~3_combout ),
	.cin(gnd),
	.combout(\Decoder0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~4 .lut_mask = 16'h4400;
defparam \Decoder0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N17
dffeas \regs[21][1] (
	.clk(CLK),
	.d(\regs[21][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][1] .is_wysiwyg = "true";
defparam \regs[21][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N18
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[21][1]~q ))) # (!dcifimemload_23 & (\regs[17][1]~q ))))

	.dataa(\regs[17][1]~q ),
	.datab(\regs[21][1]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hFC0A;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N0
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (dcifimemload_24 & ((\Mux30~0_combout  & (\regs[29][1]~q )) # (!\Mux30~0_combout  & ((\regs[25][1]~q ))))) # (!dcifimemload_24 & (((\Mux30~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[29][1]~q ),
	.datac(\regs[25][1]~q ),
	.datad(\Mux30~0_combout ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hDDA0;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N25
dffeas \regs[18][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][1] .is_wysiwyg = "true";
defparam \regs[18][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N4
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[26][1]~q )) # (!dcifimemload_24 & ((\regs[18][1]~q )))))

	.dataa(\regs[26][1]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[18][1]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hEE30;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N20
cycloneive_lcell_comb \regs[22][1]~feeder (
// Equation(s):
// \regs[22][1]~feeder_combout  = \regs~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[22][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][1]~feeder .lut_mask = 16'hF0F0;
defparam \regs[22][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \Decoder0~8 (
// Equation(s):
// \Decoder0~8_combout  = (\Selector64~0_combout  & (!\Selector65~0_combout  & (\Selector66~0_combout  & \Decoder0~7_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\Decoder0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~8 .lut_mask = 16'h2000;
defparam \Decoder0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N21
dffeas \regs[22][1] (
	.clk(CLK),
	.d(\regs[22][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][1] .is_wysiwyg = "true";
defparam \regs[22][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N6
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (dcifimemload_23 & ((\Mux30~2_combout  & (\regs[30][1]~q )) # (!\Mux30~2_combout  & ((\regs[22][1]~q ))))) # (!dcifimemload_23 & (((\Mux30~2_combout ))))

	.dataa(\regs[30][1]~q ),
	.datab(dcifimemload_23),
	.datac(\Mux30~2_combout ),
	.datad(\regs[22][1]~q ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hBCB0;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y37_N23
dffeas \regs[28][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][1] .is_wysiwyg = "true";
defparam \regs[28][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N7
dffeas \regs[20][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][1] .is_wysiwyg = "true";
defparam \regs[20][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N5
dffeas \regs[24][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][1] .is_wysiwyg = "true";
defparam \regs[24][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N4
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (dcifimemload_24 & (((\regs[24][1]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[16][1]~q  & ((!dcifimemload_23))))

	.dataa(\regs[16][1]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[24][1]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hCCE2;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N6
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// \Mux30~5_combout  = (dcifimemload_23 & ((\Mux30~4_combout  & (\regs[28][1]~q )) # (!\Mux30~4_combout  & ((\regs[20][1]~q ))))) # (!dcifimemload_23 & (((\Mux30~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[28][1]~q ),
	.datac(\regs[20][1]~q ),
	.datad(\Mux30~4_combout ),
	.cin(gnd),
	.combout(\Mux30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'hDDA0;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N28
cycloneive_lcell_comb \Mux30~6 (
// Equation(s):
// \Mux30~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux30~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux30~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux30~3_combout ),
	.datad(\Mux30~5_combout ),
	.cin(gnd),
	.combout(\Mux30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~6 .lut_mask = 16'hB9A8;
defparam \Mux30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N30
cycloneive_lcell_comb \Mux30~9 (
// Equation(s):
// \Mux30~9_combout  = (dcifimemload_21 & ((\Mux30~6_combout  & (\Mux30~8_combout )) # (!\Mux30~6_combout  & ((\Mux30~1_combout ))))) # (!dcifimemload_21 & (((\Mux30~6_combout ))))

	.dataa(\Mux30~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux30~1_combout ),
	.datad(\Mux30~6_combout ),
	.cin(gnd),
	.combout(\Mux30~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~9 .lut_mask = 16'hBBC0;
defparam \Mux30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N29
dffeas \regs[9][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][1] .is_wysiwyg = "true";
defparam \regs[9][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N15
dffeas \regs[10][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][1] .is_wysiwyg = "true";
defparam \regs[10][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N14
cycloneive_lcell_comb \Mux30~10 (
// Equation(s):
// \Mux30~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][1]~q ))) # (!dcifimemload_22 & (\regs[8][1]~q ))))

	.dataa(\regs[8][1]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[10][1]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~10 .lut_mask = 16'hFC22;
defparam \Mux30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N6
cycloneive_lcell_comb \Mux30~11 (
// Equation(s):
// \Mux30~11_combout  = (dcifimemload_21 & ((\Mux30~10_combout  & (\regs[11][1]~q )) # (!\Mux30~10_combout  & ((\regs[9][1]~q ))))) # (!dcifimemload_21 & (((\Mux30~10_combout ))))

	.dataa(\regs[11][1]~q ),
	.datab(\regs[9][1]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux30~10_combout ),
	.cin(gnd),
	.combout(\Mux30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~11 .lut_mask = 16'hAFC0;
defparam \Mux30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y31_N19
dffeas \regs[15][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][1] .is_wysiwyg = "true";
defparam \regs[15][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N29
dffeas \regs[14][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][1] .is_wysiwyg = "true";
defparam \regs[14][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N25
dffeas \regs[12][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][1] .is_wysiwyg = "true";
defparam \regs[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N2
cycloneive_lcell_comb \Decoder0~35 (
// Equation(s):
// \Decoder0~35_combout  = (!\Selector64~0_combout  & (\Selector65~0_combout  & \Decoder0~3_combout ))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(gnd),
	.datad(\Decoder0~3_combout ),
	.cin(gnd),
	.combout(\Decoder0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~35 .lut_mask = 16'h4400;
defparam \Decoder0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N7
dffeas \regs[13][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][1] .is_wysiwyg = "true";
defparam \regs[13][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N6
cycloneive_lcell_comb \Mux30~17 (
// Equation(s):
// \Mux30~17_combout  = (dcifimemload_21 & (((\regs[13][1]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][1]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][1]~q ),
	.datac(\regs[13][1]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux30~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~17 .lut_mask = 16'hAAE4;
defparam \Mux30~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N28
cycloneive_lcell_comb \Mux30~18 (
// Equation(s):
// \Mux30~18_combout  = (dcifimemload_22 & ((\Mux30~17_combout  & (\regs[15][1]~q )) # (!\Mux30~17_combout  & ((\regs[14][1]~q ))))) # (!dcifimemload_22 & (((\Mux30~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][1]~q ),
	.datac(\regs[14][1]~q ),
	.datad(\Mux30~17_combout ),
	.cin(gnd),
	.combout(\Mux30~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~18 .lut_mask = 16'hDDA0;
defparam \Mux30~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N17
dffeas \regs[3][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][1] .is_wysiwyg = "true";
defparam \regs[3][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N2
cycloneive_lcell_comb \Mux30~14 (
// Equation(s):
// \Mux30~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][1]~q ))) # (!dcifimemload_22 & (\regs[1][1]~q ))))

	.dataa(\regs[1][1]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[3][1]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux30~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~14 .lut_mask = 16'hC088;
defparam \Mux30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N26
cycloneive_lcell_comb \Mux30~15 (
// Equation(s):
// \Mux30~15_combout  = (\Mux30~14_combout ) # ((\regs[2][1]~q  & (!dcifimemload_21 & dcifimemload_22)))

	.dataa(\regs[2][1]~q ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\Mux30~14_combout ),
	.cin(gnd),
	.combout(\Mux30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~15 .lut_mask = 16'hFF20;
defparam \Mux30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N15
dffeas \regs[7][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][1] .is_wysiwyg = "true";
defparam \regs[7][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \Decoder0~27 (
// Equation(s):
// \Decoder0~27_combout  = (!\Selector64~0_combout  & (!\Selector65~0_combout  & (\Selector66~0_combout  & \Decoder0~7_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\Decoder0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~27 .lut_mask = 16'h1000;
defparam \Decoder0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N13
dffeas \regs[6][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][1] .is_wysiwyg = "true";
defparam \regs[6][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N13
dffeas \regs[5][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][1] .is_wysiwyg = "true";
defparam \regs[5][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \Mux30~12 (
// Equation(s):
// \Mux30~12_combout  = (dcifimemload_21 & (((\regs[5][1]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][1]~q  & ((!dcifimemload_22))))

	.dataa(\regs[4][1]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[5][1]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~12 .lut_mask = 16'hCCE2;
defparam \Mux30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N12
cycloneive_lcell_comb \Mux30~13 (
// Equation(s):
// \Mux30~13_combout  = (dcifimemload_22 & ((\Mux30~12_combout  & (\regs[7][1]~q )) # (!\Mux30~12_combout  & ((\regs[6][1]~q ))))) # (!dcifimemload_22 & (((\Mux30~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[7][1]~q ),
	.datac(\regs[6][1]~q ),
	.datad(\Mux30~12_combout ),
	.cin(gnd),
	.combout(\Mux30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~13 .lut_mask = 16'hDDA0;
defparam \Mux30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N20
cycloneive_lcell_comb \Mux30~16 (
// Equation(s):
// \Mux30~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux30~13_combout ))) # (!dcifimemload_23 & (\Mux30~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux30~15_combout ),
	.datad(\Mux30~13_combout ),
	.cin(gnd),
	.combout(\Mux30~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~16 .lut_mask = 16'hDC98;
defparam \Mux30~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N6
cycloneive_lcell_comb \Mux30~19 (
// Equation(s):
// \Mux30~19_combout  = (dcifimemload_24 & ((\Mux30~16_combout  & ((\Mux30~18_combout ))) # (!\Mux30~16_combout  & (\Mux30~11_combout )))) # (!dcifimemload_24 & (((\Mux30~16_combout ))))

	.dataa(\Mux30~11_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux30~18_combout ),
	.datad(\Mux30~16_combout ),
	.cin(gnd),
	.combout(\Mux30~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~19 .lut_mask = 16'hF388;
defparam \Mux30~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N14
cycloneive_lcell_comb \regs~8 (
// Equation(s):
// \regs~8_combout  = (!\Equal0~1_combout  & \Selector1~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Equal0~1_combout ),
	.datad(Selector1),
	.cin(gnd),
	.combout(\regs~8_combout ),
	.cout());
// synopsys translate_off
defparam \regs~8 .lut_mask = 16'h0F00;
defparam \regs~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N3
dffeas \regs[31][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][30] .is_wysiwyg = "true";
defparam \regs[31][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N23
dffeas \regs[27][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][30] .is_wysiwyg = "true";
defparam \regs[27][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N25
dffeas \regs[23][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][30] .is_wysiwyg = "true";
defparam \regs[23][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N24
cycloneive_lcell_comb \Mux33~7 (
// Equation(s):
// \Mux33~7_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\regs[23][30]~q ))) # (!dcifimemload_18 & (\regs[19][30]~q ))))

	.dataa(\regs[19][30]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[23][30]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux33~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~7 .lut_mask = 16'hFC22;
defparam \Mux33~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N22
cycloneive_lcell_comb \Mux33~8 (
// Equation(s):
// \Mux33~8_combout  = (dcifimemload_19 & ((\Mux33~7_combout  & (\regs[31][30]~q )) # (!\Mux33~7_combout  & ((\regs[27][30]~q ))))) # (!dcifimemload_19 & (((\Mux33~7_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[31][30]~q ),
	.datac(\regs[27][30]~q ),
	.datad(\Mux33~7_combout ),
	.cin(gnd),
	.combout(\Mux33~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~8 .lut_mask = 16'hDDA0;
defparam \Mux33~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N1
dffeas \regs[21][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][30] .is_wysiwyg = "true";
defparam \regs[21][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N0
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (dcifimemload_18 & (((\regs[21][30]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[17][30]~q  & ((!dcifimemload_19))))

	.dataa(\regs[17][30]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[21][30]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hCCE2;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N29
dffeas \regs[29][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][30] .is_wysiwyg = "true";
defparam \regs[29][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N9
dffeas \regs[25][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][30] .is_wysiwyg = "true";
defparam \regs[25][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N8
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (\Mux33~0_combout  & ((\regs[29][30]~q ) # ((!dcifimemload_19)))) # (!\Mux33~0_combout  & (((\regs[25][30]~q  & dcifimemload_19))))

	.dataa(\Mux33~0_combout ),
	.datab(\regs[29][30]~q ),
	.datac(\regs[25][30]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hD8AA;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N17
dffeas \regs[16][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][30] .is_wysiwyg = "true";
defparam \regs[16][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N15
dffeas \regs[24][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][30] .is_wysiwyg = "true";
defparam \regs[24][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N14
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[24][30]~q ))) # (!dcifimemload_19 & (\regs[16][30]~q ))))

	.dataa(dcifimemload_18),
	.datab(\regs[16][30]~q ),
	.datac(\regs[24][30]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'hFA44;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N9
dffeas \regs[20][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][30] .is_wysiwyg = "true";
defparam \regs[20][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y42_N7
dffeas \regs[28][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][30] .is_wysiwyg = "true";
defparam \regs[28][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N8
cycloneive_lcell_comb \Mux33~5 (
// Equation(s):
// \Mux33~5_combout  = (dcifimemload_18 & ((\Mux33~4_combout  & ((\regs[28][30]~q ))) # (!\Mux33~4_combout  & (\regs[20][30]~q )))) # (!dcifimemload_18 & (\Mux33~4_combout ))

	.dataa(dcifimemload_18),
	.datab(\Mux33~4_combout ),
	.datac(\regs[20][30]~q ),
	.datad(\regs[28][30]~q ),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~5 .lut_mask = 16'hEC64;
defparam \Mux33~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N2
cycloneive_lcell_comb \regs[22][30]~feeder (
// Equation(s):
// \regs[22][30]~feeder_combout  = \regs~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[22][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][30]~feeder .lut_mask = 16'hF0F0;
defparam \regs[22][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y43_N3
dffeas \regs[22][30] (
	.clk(CLK),
	.d(\regs[22][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][30] .is_wysiwyg = "true";
defparam \regs[22][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N20
cycloneive_lcell_comb \Decoder0~9 (
// Equation(s):
// \Decoder0~9_combout  = (\Selector64~0_combout  & (!\Selector66~0_combout  & (\Selector65~0_combout  & \Decoder0~7_combout )))

	.dataa(Selector64),
	.datab(Selector66),
	.datac(Selector65),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\Decoder0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~9 .lut_mask = 16'h2000;
defparam \Decoder0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y43_N29
dffeas \regs[26][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][30] .is_wysiwyg = "true";
defparam \regs[26][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N28
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[26][30]~q ))) # (!dcifimemload_19 & (\regs[18][30]~q ))))

	.dataa(\regs[18][30]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[26][30]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hFC22;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N28
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (dcifimemload_18 & ((\Mux33~2_combout  & (\regs[30][30]~q )) # (!\Mux33~2_combout  & ((\regs[22][30]~q ))))) # (!dcifimemload_18 & (((\Mux33~2_combout ))))

	.dataa(\regs[30][30]~q ),
	.datab(\regs[22][30]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux33~2_combout ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hAFC0;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N24
cycloneive_lcell_comb \Mux33~6 (
// Equation(s):
// \Mux33~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux33~3_combout ))) # (!dcifimemload_17 & (\Mux33~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux33~5_combout ),
	.datad(\Mux33~3_combout ),
	.cin(gnd),
	.combout(\Mux33~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~6 .lut_mask = 16'hDC98;
defparam \Mux33~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N5
dffeas \regs[14][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][30] .is_wysiwyg = "true";
defparam \regs[14][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N31
dffeas \regs[15][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][30] .is_wysiwyg = "true";
defparam \regs[15][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N3
dffeas \regs[13][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][30] .is_wysiwyg = "true";
defparam \regs[13][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N21
dffeas \regs[12][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][30] .is_wysiwyg = "true";
defparam \regs[12][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N20
cycloneive_lcell_comb \Mux33~17 (
// Equation(s):
// \Mux33~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][30]~q )) # (!dcifimemload_16 & ((\regs[12][30]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[13][30]~q ),
	.datac(\regs[12][30]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux33~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~17 .lut_mask = 16'hEE50;
defparam \Mux33~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N30
cycloneive_lcell_comb \Mux33~18 (
// Equation(s):
// \Mux33~18_combout  = (dcifimemload_17 & ((\Mux33~17_combout  & ((\regs[15][30]~q ))) # (!\Mux33~17_combout  & (\regs[14][30]~q )))) # (!dcifimemload_17 & (((\Mux33~17_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[14][30]~q ),
	.datac(\regs[15][30]~q ),
	.datad(\Mux33~17_combout ),
	.cin(gnd),
	.combout(\Mux33~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~18 .lut_mask = 16'hF588;
defparam \Mux33~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N11
dffeas \regs[10][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][30] .is_wysiwyg = "true";
defparam \regs[10][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N10
cycloneive_lcell_comb \Mux33~10 (
// Equation(s):
// \Mux33~10_combout  = (dcifimemload_17 & (((\regs[10][30]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\regs[8][30]~q  & ((!dcifimemload_16))))

	.dataa(\regs[8][30]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[10][30]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux33~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~10 .lut_mask = 16'hCCE2;
defparam \Mux33~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N10
cycloneive_lcell_comb \regs[11][30]~feeder (
// Equation(s):
// \regs[11][30]~feeder_combout  = \regs~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[11][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][30]~feeder .lut_mask = 16'hF0F0;
defparam \regs[11][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N11
dffeas \regs[11][30] (
	.clk(CLK),
	.d(\regs[11][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][30] .is_wysiwyg = "true";
defparam \regs[11][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N1
dffeas \regs[9][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][30] .is_wysiwyg = "true";
defparam \regs[9][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N0
cycloneive_lcell_comb \Mux33~11 (
// Equation(s):
// \Mux33~11_combout  = (\Mux33~10_combout  & ((\regs[11][30]~q ) # ((!dcifimemload_16)))) # (!\Mux33~10_combout  & (((\regs[9][30]~q  & dcifimemload_16))))

	.dataa(\Mux33~10_combout ),
	.datab(\regs[11][30]~q ),
	.datac(\regs[9][30]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux33~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~11 .lut_mask = 16'hD8AA;
defparam \Mux33~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N29
dffeas \regs[6][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][30] .is_wysiwyg = "true";
defparam \regs[6][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N31
dffeas \regs[7][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][30] .is_wysiwyg = "true";
defparam \regs[7][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N21
dffeas \regs[4][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][30] .is_wysiwyg = "true";
defparam \regs[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N20
cycloneive_lcell_comb \Mux33~12 (
// Equation(s):
// \Mux33~12_combout  = (dcifimemload_16 & ((\regs[5][30]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][30]~q  & !dcifimemload_17))))

	.dataa(\regs[5][30]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][30]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux33~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~12 .lut_mask = 16'hCCB8;
defparam \Mux33~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N30
cycloneive_lcell_comb \Mux33~13 (
// Equation(s):
// \Mux33~13_combout  = (dcifimemload_17 & ((\Mux33~12_combout  & ((\regs[7][30]~q ))) # (!\Mux33~12_combout  & (\regs[6][30]~q )))) # (!dcifimemload_17 & (((\Mux33~12_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][30]~q ),
	.datac(\regs[7][30]~q ),
	.datad(\Mux33~12_combout ),
	.cin(gnd),
	.combout(\Mux33~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~13 .lut_mask = 16'hF588;
defparam \Mux33~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N14
cycloneive_lcell_comb \Decoder0~32 (
// Equation(s):
// \Decoder0~32_combout  = (!\Selector64~0_combout  & (!\Selector65~0_combout  & (!\Selector66~0_combout  & \Decoder0~7_combout )))

	.dataa(Selector64),
	.datab(Selector65),
	.datac(Selector66),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\Decoder0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~32 .lut_mask = 16'h0100;
defparam \Decoder0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N19
dffeas \regs[2][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][30] .is_wysiwyg = "true";
defparam \regs[2][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N28
cycloneive_lcell_comb \regs[3][30]~feeder (
// Equation(s):
// \regs[3][30]~feeder_combout  = \regs~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[3][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][30]~feeder .lut_mask = 16'hF0F0;
defparam \regs[3][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N29
dffeas \regs[3][30] (
	.clk(CLK),
	.d(\regs[3][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][30] .is_wysiwyg = "true";
defparam \regs[3][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N1
dffeas \regs[1][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][30] .is_wysiwyg = "true";
defparam \regs[1][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N0
cycloneive_lcell_comb \Mux33~14 (
// Equation(s):
// \Mux33~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][30]~q )) # (!dcifimemload_17 & ((\regs[1][30]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[3][30]~q ),
	.datac(\regs[1][30]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux33~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~14 .lut_mask = 16'hD800;
defparam \Mux33~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N18
cycloneive_lcell_comb \Mux33~15 (
// Equation(s):
// \Mux33~15_combout  = (\Mux33~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][30]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][30]~q ),
	.datad(\Mux33~14_combout ),
	.cin(gnd),
	.combout(\Mux33~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~15 .lut_mask = 16'hFF40;
defparam \Mux33~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N20
cycloneive_lcell_comb \Mux33~16 (
// Equation(s):
// \Mux33~16_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\Mux33~13_combout )) # (!dcifimemload_18 & ((\Mux33~15_combout )))))

	.dataa(\Mux33~13_combout ),
	.datab(dcifimemload_19),
	.datac(dcifimemload_18),
	.datad(\Mux33~15_combout ),
	.cin(gnd),
	.combout(\Mux33~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~16 .lut_mask = 16'hE3E0;
defparam \Mux33~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N2
cycloneive_lcell_comb \Mux1~14 (
// Equation(s):
// \Mux1~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][30]~q ))) # (!dcifimemload_22 & (\regs[1][30]~q ))))

	.dataa(\regs[1][30]~q ),
	.datab(\regs[3][30]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~14 .lut_mask = 16'hC0A0;
defparam \Mux1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N4
cycloneive_lcell_comb \Mux1~15 (
// Equation(s):
// \Mux1~15_combout  = (\Mux1~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][30]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux1~14_combout ),
	.datad(\regs[2][30]~q ),
	.cin(gnd),
	.combout(\Mux1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~15 .lut_mask = 16'hF2F0;
defparam \Mux1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N28
cycloneive_lcell_comb \regs[8][30]~feeder (
// Equation(s):
// \regs[8][30]~feeder_combout  = \regs~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~8_combout ),
	.cin(gnd),
	.combout(\regs[8][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][30]~feeder .lut_mask = 16'hFF00;
defparam \regs[8][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y42_N29
dffeas \regs[8][30] (
	.clk(CLK),
	.d(\regs[8][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][30] .is_wysiwyg = "true";
defparam \regs[8][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N16
cycloneive_lcell_comb \Mux1~12 (
// Equation(s):
// \Mux1~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\regs[10][30]~q )) # (!dcifimemload_22 & ((\regs[8][30]~q )))))

	.dataa(\regs[10][30]~q ),
	.datab(\regs[8][30]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~12 .lut_mask = 16'hFA0C;
defparam \Mux1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N18
cycloneive_lcell_comb \Mux1~13 (
// Equation(s):
// \Mux1~13_combout  = (dcifimemload_21 & ((\Mux1~12_combout  & (\regs[11][30]~q )) # (!\Mux1~12_combout  & ((\regs[9][30]~q ))))) # (!dcifimemload_21 & (((\Mux1~12_combout ))))

	.dataa(\regs[11][30]~q ),
	.datab(\regs[9][30]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux1~12_combout ),
	.cin(gnd),
	.combout(\Mux1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~13 .lut_mask = 16'hAFC0;
defparam \Mux1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N14
cycloneive_lcell_comb \Mux1~16 (
// Equation(s):
// \Mux1~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux1~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & (\Mux1~15_combout )))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux1~15_combout ),
	.datad(\Mux1~13_combout ),
	.cin(gnd),
	.combout(\Mux1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~16 .lut_mask = 16'hBA98;
defparam \Mux1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N2
cycloneive_lcell_comb \Mux1~17 (
// Equation(s):
// \Mux1~17_combout  = (dcifimemload_21 & (((\regs[13][30]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][30]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][30]~q ),
	.datac(\regs[13][30]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~17 .lut_mask = 16'hAAE4;
defparam \Mux1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N4
cycloneive_lcell_comb \Mux1~18 (
// Equation(s):
// \Mux1~18_combout  = (dcifimemload_22 & ((\Mux1~17_combout  & (\regs[15][30]~q )) # (!\Mux1~17_combout  & ((\regs[14][30]~q ))))) # (!dcifimemload_22 & (((\Mux1~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][30]~q ),
	.datac(\regs[14][30]~q ),
	.datad(\Mux1~17_combout ),
	.cin(gnd),
	.combout(\Mux1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~18 .lut_mask = 16'hDDA0;
defparam \Mux1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N11
dffeas \regs[5][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][30] .is_wysiwyg = "true";
defparam \regs[5][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N10
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// \Mux1~10_combout  = (dcifimemload_21 & (((\regs[5][30]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][30]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][30]~q ),
	.datac(\regs[5][30]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hAAE4;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N28
cycloneive_lcell_comb \Mux1~11 (
// Equation(s):
// \Mux1~11_combout  = (dcifimemload_22 & ((\Mux1~10_combout  & (\regs[7][30]~q )) # (!\Mux1~10_combout  & ((\regs[6][30]~q ))))) # (!dcifimemload_22 & (((\Mux1~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[7][30]~q ),
	.datac(\regs[6][30]~q ),
	.datad(\Mux1~10_combout ),
	.cin(gnd),
	.combout(\Mux1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~11 .lut_mask = 16'hDDA0;
defparam \Mux1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N8
cycloneive_lcell_comb \Mux1~19 (
// Equation(s):
// \Mux1~19_combout  = (dcifimemload_23 & ((\Mux1~16_combout  & (\Mux1~18_combout )) # (!\Mux1~16_combout  & ((\Mux1~11_combout ))))) # (!dcifimemload_23 & (\Mux1~16_combout ))

	.dataa(dcifimemload_23),
	.datab(\Mux1~16_combout ),
	.datac(\Mux1~18_combout ),
	.datad(\Mux1~11_combout ),
	.cin(gnd),
	.combout(\Mux1~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~19 .lut_mask = 16'hE6C4;
defparam \Mux1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N8
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (dcifimemload_24 & (((\regs[25][30]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[17][30]~q  & ((!dcifimemload_23))))

	.dataa(\regs[17][30]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[25][30]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hCCE2;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N28
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (dcifimemload_23 & ((\Mux1~0_combout  & ((\regs[29][30]~q ))) # (!\Mux1~0_combout  & (\regs[21][30]~q )))) # (!dcifimemload_23 & (((\Mux1~0_combout ))))

	.dataa(\regs[21][30]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[29][30]~q ),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hF388;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N9
dffeas \regs[19][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][30] .is_wysiwyg = "true";
defparam \regs[19][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N8
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (dcifimemload_24 & ((\regs[27][30]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[19][30]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][30]~q ),
	.datac(\regs[19][30]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hAAD8;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N2
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (\Mux1~7_combout  & (((\regs[31][30]~q ) # (!dcifimemload_23)))) # (!\Mux1~7_combout  & (\regs[23][30]~q  & ((dcifimemload_23))))

	.dataa(\regs[23][30]~q ),
	.datab(\Mux1~7_combout ),
	.datac(\regs[31][30]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hE2CC;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N28
cycloneive_lcell_comb \regs[30][30]~feeder (
// Equation(s):
// \regs[30][30]~feeder_combout  = \regs~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~8_combout ),
	.cin(gnd),
	.combout(\regs[30][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[30][30]~feeder .lut_mask = 16'hFF00;
defparam \regs[30][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y43_N29
dffeas \regs[30][30] (
	.clk(CLK),
	.d(\regs[30][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][30] .is_wysiwyg = "true";
defparam \regs[30][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N22
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (dcifimemload_23 & (((\regs[22][30]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[18][30]~q  & ((!dcifimemload_24))))

	.dataa(\regs[18][30]~q ),
	.datab(\regs[22][30]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hF0CA;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N18
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (dcifimemload_24 & ((\Mux1~2_combout  & ((\regs[30][30]~q ))) # (!\Mux1~2_combout  & (\regs[26][30]~q )))) # (!dcifimemload_24 & (((\Mux1~2_combout ))))

	.dataa(\regs[26][30]~q ),
	.datab(\regs[30][30]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux1~2_combout ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hCFA0;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N16
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (dcifimemload_23 & ((\regs[20][30]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[16][30]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[20][30]~q ),
	.datac(\regs[16][30]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hAAD8;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N6
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (dcifimemload_24 & ((\Mux1~4_combout  & ((\regs[28][30]~q ))) # (!\Mux1~4_combout  & (\regs[24][30]~q )))) # (!dcifimemload_24 & (((\Mux1~4_combout ))))

	.dataa(\regs[24][30]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[28][30]~q ),
	.datad(\Mux1~4_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hF388;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N24
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux1~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux1~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux1~3_combout ),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hB9A8;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N10
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// \Mux1~9_combout  = (dcifimemload_21 & ((\Mux1~6_combout  & ((\Mux1~8_combout ))) # (!\Mux1~6_combout  & (\Mux1~1_combout )))) # (!dcifimemload_21 & (((\Mux1~6_combout ))))

	.dataa(\Mux1~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux1~8_combout ),
	.datad(\Mux1~6_combout ),
	.cin(gnd),
	.combout(\Mux1~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hF388;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N0
cycloneive_lcell_comb \regs~9 (
// Equation(s):
// \regs~9_combout  = (!\Equal0~1_combout  & \Selector2~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Equal0~1_combout ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\regs~9_combout ),
	.cout());
// synopsys translate_off
defparam \regs~9 .lut_mask = 16'h0F00;
defparam \regs~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N27
dffeas \regs[31][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][29] .is_wysiwyg = "true";
defparam \regs[31][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N8
cycloneive_lcell_comb \regs[23][29]~feeder (
// Equation(s):
// \regs[23][29]~feeder_combout  = \regs~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~9_combout ),
	.cin(gnd),
	.combout(\regs[23][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][29]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N9
dffeas \regs[23][29] (
	.clk(CLK),
	.d(\regs[23][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][29] .is_wysiwyg = "true";
defparam \regs[23][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N2
cycloneive_lcell_comb \regs[27][29]~feeder (
// Equation(s):
// \regs[27][29]~feeder_combout  = \regs~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~9_combout ),
	.cin(gnd),
	.combout(\regs[27][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][29]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N3
dffeas \regs[27][29] (
	.clk(CLK),
	.d(\regs[27][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][29] .is_wysiwyg = "true";
defparam \regs[27][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N24
cycloneive_lcell_comb \Mux34~7 (
// Equation(s):
// \Mux34~7_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[27][29]~q ))) # (!dcifimemload_19 & (\regs[19][29]~q ))))

	.dataa(\regs[19][29]~q ),
	.datab(\regs[27][29]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux34~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~7 .lut_mask = 16'hFC0A;
defparam \Mux34~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N26
cycloneive_lcell_comb \Mux34~8 (
// Equation(s):
// \Mux34~8_combout  = (dcifimemload_18 & ((\Mux34~7_combout  & (\regs[31][29]~q )) # (!\Mux34~7_combout  & ((\regs[23][29]~q ))))) # (!dcifimemload_18 & (((\Mux34~7_combout ))))

	.dataa(\regs[31][29]~q ),
	.datab(\regs[23][29]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux34~7_combout ),
	.cin(gnd),
	.combout(\Mux34~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~8 .lut_mask = 16'hAFC0;
defparam \Mux34~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N18
cycloneive_lcell_comb \regs[21][29]~feeder (
// Equation(s):
// \regs[21][29]~feeder_combout  = \regs~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[21][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][29]~feeder .lut_mask = 16'hF0F0;
defparam \regs[21][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N19
dffeas \regs[21][29] (
	.clk(CLK),
	.d(\regs[21][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][29] .is_wysiwyg = "true";
defparam \regs[21][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N25
dffeas \regs[25][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][29] .is_wysiwyg = "true";
defparam \regs[25][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N24
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[25][29]~q ))) # (!dcifimemload_19 & (\regs[17][29]~q ))))

	.dataa(\regs[17][29]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[25][29]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hFC22;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N1
dffeas \regs[29][29] (
	.clk(CLK),
	.d(\regs~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][29] .is_wysiwyg = "true";
defparam \regs[29][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N20
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (dcifimemload_18 & ((\Mux34~0_combout  & ((\regs[29][29]~q ))) # (!\Mux34~0_combout  & (\regs[21][29]~q )))) # (!dcifimemload_18 & (((\Mux34~0_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[21][29]~q ),
	.datac(\Mux34~0_combout ),
	.datad(\regs[29][29]~q ),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hF858;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N15
dffeas \regs[28][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][29] .is_wysiwyg = "true";
defparam \regs[28][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N31
dffeas \regs[24][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][29] .is_wysiwyg = "true";
defparam \regs[24][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N13
dffeas \regs[20][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][29] .is_wysiwyg = "true";
defparam \regs[20][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N12
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (dcifimemload_18 & (((\regs[20][29]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[16][29]~q  & ((!dcifimemload_19))))

	.dataa(\regs[16][29]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[20][29]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'hCCE2;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N30
cycloneive_lcell_comb \Mux34~5 (
// Equation(s):
// \Mux34~5_combout  = (dcifimemload_19 & ((\Mux34~4_combout  & (\regs[28][29]~q )) # (!\Mux34~4_combout  & ((\regs[24][29]~q ))))) # (!dcifimemload_19 & (((\Mux34~4_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[28][29]~q ),
	.datac(\regs[24][29]~q ),
	.datad(\Mux34~4_combout ),
	.cin(gnd),
	.combout(\Mux34~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~5 .lut_mask = 16'hDDA0;
defparam \Mux34~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N27
dffeas \regs[30][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][29] .is_wysiwyg = "true";
defparam \regs[30][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y43_N17
dffeas \regs[22][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][29] .is_wysiwyg = "true";
defparam \regs[22][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N16
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (dcifimemload_18 & (((\regs[22][29]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[18][29]~q  & ((!dcifimemload_19))))

	.dataa(\regs[18][29]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[22][29]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hCCE2;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N2
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (dcifimemload_19 & ((\Mux34~2_combout  & ((\regs[30][29]~q ))) # (!\Mux34~2_combout  & (\regs[26][29]~q )))) # (!dcifimemload_19 & (((\Mux34~2_combout ))))

	.dataa(\regs[26][29]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[30][29]~q ),
	.datad(\Mux34~2_combout ),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hF388;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N10
cycloneive_lcell_comb \Mux34~6 (
// Equation(s):
// \Mux34~6_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux34~3_combout ))) # (!dcifimemload_17 & (\Mux34~5_combout ))))

	.dataa(\Mux34~5_combout ),
	.datab(dcifimemload_16),
	.datac(dcifimemload_17),
	.datad(\Mux34~3_combout ),
	.cin(gnd),
	.combout(\Mux34~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~6 .lut_mask = 16'hF2C2;
defparam \Mux34~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N23
dffeas \regs[5][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][29] .is_wysiwyg = "true";
defparam \regs[5][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N22
cycloneive_lcell_comb \Mux34~10 (
// Equation(s):
// \Mux34~10_combout  = (dcifimemload_16 & (((\regs[5][29]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][29]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][29]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[5][29]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux34~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~10 .lut_mask = 16'hCCE2;
defparam \Mux34~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N15
dffeas \regs[7][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][29] .is_wysiwyg = "true";
defparam \regs[7][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N5
dffeas \regs[6][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][29] .is_wysiwyg = "true";
defparam \regs[6][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N4
cycloneive_lcell_comb \Mux34~11 (
// Equation(s):
// \Mux34~11_combout  = (\Mux34~10_combout  & ((\regs[7][29]~q ) # ((!dcifimemload_17)))) # (!\Mux34~10_combout  & (((\regs[6][29]~q  & dcifimemload_17))))

	.dataa(\Mux34~10_combout ),
	.datab(\regs[7][29]~q ),
	.datac(\regs[6][29]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux34~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~11 .lut_mask = 16'hD8AA;
defparam \Mux34~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N13
dffeas \regs[14][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][29] .is_wysiwyg = "true";
defparam \regs[14][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N19
dffeas \regs[13][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][29] .is_wysiwyg = "true";
defparam \regs[13][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N9
dffeas \regs[12][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][29] .is_wysiwyg = "true";
defparam \regs[12][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N8
cycloneive_lcell_comb \Mux34~17 (
// Equation(s):
// \Mux34~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][29]~q )) # (!dcifimemload_16 & ((\regs[12][29]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[13][29]~q ),
	.datac(\regs[12][29]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux34~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~17 .lut_mask = 16'hEE50;
defparam \Mux34~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y31_N23
dffeas \regs[15][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][29] .is_wysiwyg = "true";
defparam \regs[15][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N22
cycloneive_lcell_comb \Mux34~18 (
// Equation(s):
// \Mux34~18_combout  = (\Mux34~17_combout  & (((\regs[15][29]~q ) # (!dcifimemload_17)))) # (!\Mux34~17_combout  & (\regs[14][29]~q  & ((dcifimemload_17))))

	.dataa(\regs[14][29]~q ),
	.datab(\Mux34~17_combout ),
	.datac(\regs[15][29]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux34~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~18 .lut_mask = 16'hE2CC;
defparam \Mux34~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N13
dffeas \regs[3][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][29] .is_wysiwyg = "true";
defparam \regs[3][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N15
dffeas \regs[1][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][29] .is_wysiwyg = "true";
defparam \regs[1][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N14
cycloneive_lcell_comb \Mux34~14 (
// Equation(s):
// \Mux34~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][29]~q )) # (!dcifimemload_17 & ((\regs[1][29]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[3][29]~q ),
	.datac(\regs[1][29]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux34~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~14 .lut_mask = 16'hD800;
defparam \Mux34~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N21
dffeas \regs[2][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][29] .is_wysiwyg = "true";
defparam \regs[2][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N20
cycloneive_lcell_comb \Mux34~15 (
// Equation(s):
// \Mux34~15_combout  = (\Mux34~14_combout ) # ((dcifimemload_17 & (\regs[2][29]~q  & !dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\Mux34~14_combout ),
	.datac(\regs[2][29]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux34~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~15 .lut_mask = 16'hCCEC;
defparam \Mux34~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N9
dffeas \regs[9][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][29] .is_wysiwyg = "true";
defparam \regs[9][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N11
dffeas \regs[11][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][29] .is_wysiwyg = "true";
defparam \regs[11][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N1
dffeas \regs[8][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][29] .is_wysiwyg = "true";
defparam \regs[8][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N0
cycloneive_lcell_comb \Mux34~12 (
// Equation(s):
// \Mux34~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][29]~q )) # (!dcifimemload_17 & ((\regs[8][29]~q )))))

	.dataa(\regs[10][29]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[8][29]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux34~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~12 .lut_mask = 16'hEE30;
defparam \Mux34~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N10
cycloneive_lcell_comb \Mux34~13 (
// Equation(s):
// \Mux34~13_combout  = (dcifimemload_16 & ((\Mux34~12_combout  & ((\regs[11][29]~q ))) # (!\Mux34~12_combout  & (\regs[9][29]~q )))) # (!dcifimemload_16 & (((\Mux34~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][29]~q ),
	.datac(\regs[11][29]~q ),
	.datad(\Mux34~12_combout ),
	.cin(gnd),
	.combout(\Mux34~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~13 .lut_mask = 16'hF588;
defparam \Mux34~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N18
cycloneive_lcell_comb \Mux34~16 (
// Equation(s):
// \Mux34~16_combout  = (dcifimemload_19 & (((dcifimemload_18) # (\Mux34~13_combout )))) # (!dcifimemload_19 & (\Mux34~15_combout  & (!dcifimemload_18)))

	.dataa(\Mux34~15_combout ),
	.datab(dcifimemload_19),
	.datac(dcifimemload_18),
	.datad(\Mux34~13_combout ),
	.cin(gnd),
	.combout(\Mux34~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~16 .lut_mask = 16'hCEC2;
defparam \Mux34~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N9
dffeas \regs[16][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][29] .is_wysiwyg = "true";
defparam \regs[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N8
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[24][29]~q )) # (!dcifimemload_24 & ((\regs[16][29]~q )))))

	.dataa(\regs[24][29]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[16][29]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hEE30;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N14
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (\Mux2~4_combout  & (((\regs[28][29]~q ) # (!dcifimemload_23)))) # (!\Mux2~4_combout  & (\regs[20][29]~q  & ((dcifimemload_23))))

	.dataa(\regs[20][29]~q ),
	.datab(\Mux2~4_combout ),
	.datac(\regs[28][29]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hE2CC;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N17
dffeas \regs[18][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][29] .is_wysiwyg = "true";
defparam \regs[18][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N16
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[26][29]~q )) # (!dcifimemload_24 & ((\regs[18][29]~q )))))

	.dataa(\regs[26][29]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[18][29]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hEE30;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N26
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (dcifimemload_23 & ((\Mux2~2_combout  & ((\regs[30][29]~q ))) # (!\Mux2~2_combout  & (\regs[22][29]~q )))) # (!dcifimemload_23 & (((\Mux2~2_combout ))))

	.dataa(\regs[22][29]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[30][29]~q ),
	.datad(\Mux2~2_combout ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hF388;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N22
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux2~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux2~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux2~5_combout ),
	.datad(\Mux2~3_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hBA98;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N29
dffeas \regs[19][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][29] .is_wysiwyg = "true";
defparam \regs[19][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N28
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[23][29]~q )) # (!dcifimemload_23 & ((\regs[19][29]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[23][29]~q ),
	.datac(\regs[19][29]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hEE50;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N26
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (dcifimemload_24 & ((\Mux2~7_combout  & ((\regs[31][29]~q ))) # (!\Mux2~7_combout  & (\regs[27][29]~q )))) # (!dcifimemload_24 & (((\Mux2~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][29]~q ),
	.datac(\regs[31][29]~q ),
	.datad(\Mux2~7_combout ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hF588;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N1
dffeas \regs[17][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][29] .is_wysiwyg = "true";
defparam \regs[17][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N10
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (dcifimemload_23 & ((\regs[21][29]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[17][29]~q  & !dcifimemload_24))))

	.dataa(\regs[21][29]~q ),
	.datab(\regs[17][29]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hF0AC;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N22
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (\Mux2~0_combout  & ((\regs[29][29]~q ) # ((!dcifimemload_24)))) # (!\Mux2~0_combout  & (((\regs[25][29]~q  & dcifimemload_24))))

	.dataa(\regs[29][29]~q ),
	.datab(\regs[25][29]~q ),
	.datac(\Mux2~0_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hACF0;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N8
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// \Mux2~9_combout  = (\Mux2~6_combout  & (((\Mux2~8_combout )) # (!dcifimemload_21))) # (!\Mux2~6_combout  & (dcifimemload_21 & ((\Mux2~1_combout ))))

	.dataa(\Mux2~6_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux2~8_combout ),
	.datad(\Mux2~1_combout ),
	.cin(gnd),
	.combout(\Mux2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hE6A2;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N18
cycloneive_lcell_comb \Mux2~17 (
// Equation(s):
// \Mux2~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\regs[13][29]~q ))) # (!dcifimemload_21 & (\regs[12][29]~q ))))

	.dataa(\regs[12][29]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[13][29]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~17 .lut_mask = 16'hFC22;
defparam \Mux2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N12
cycloneive_lcell_comb \Mux2~18 (
// Equation(s):
// \Mux2~18_combout  = (dcifimemload_22 & ((\Mux2~17_combout  & (\regs[15][29]~q )) # (!\Mux2~17_combout  & ((\regs[14][29]~q ))))) # (!dcifimemload_22 & (((\Mux2~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][29]~q ),
	.datac(\regs[14][29]~q ),
	.datad(\Mux2~17_combout ),
	.cin(gnd),
	.combout(\Mux2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~18 .lut_mask = 16'hDDA0;
defparam \Mux2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N11
dffeas \regs[10][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][29] .is_wysiwyg = "true";
defparam \regs[10][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N10
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\regs[10][29]~q )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\regs[8][29]~q ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[10][29]~q ),
	.datad(\regs[8][29]~q ),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hB9A8;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N8
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (dcifimemload_21 & ((\Mux2~10_combout  & (\regs[11][29]~q )) # (!\Mux2~10_combout  & ((\regs[9][29]~q ))))) # (!dcifimemload_21 & (((\Mux2~10_combout ))))

	.dataa(\regs[11][29]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[9][29]~q ),
	.datad(\Mux2~10_combout ),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hBBC0;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N12
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// \Mux2~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][29]~q ))) # (!dcifimemload_22 & (\regs[1][29]~q ))))

	.dataa(\regs[1][29]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[3][29]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'hC088;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N26
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (\Mux2~14_combout ) # ((\regs[2][29]~q  & (!dcifimemload_21 & dcifimemload_22)))

	.dataa(\regs[2][29]~q ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\Mux2~14_combout ),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hFF20;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N5
dffeas \regs[4][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][29] .is_wysiwyg = "true";
defparam \regs[4][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N4
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (dcifimemload_21 & ((dcifimemload_22) # ((\regs[5][29]~q )))) # (!dcifimemload_21 & (!dcifimemload_22 & (\regs[4][29]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[4][29]~q ),
	.datad(\regs[5][29]~q ),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hBA98;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N14
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (dcifimemload_22 & ((\Mux2~12_combout  & ((\regs[7][29]~q ))) # (!\Mux2~12_combout  & (\regs[6][29]~q )))) # (!dcifimemload_22 & (((\Mux2~12_combout ))))

	.dataa(\regs[6][29]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[7][29]~q ),
	.datad(\Mux2~12_combout ),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hF388;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N10
cycloneive_lcell_comb \Mux2~16 (
// Equation(s):
// \Mux2~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux2~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & (\Mux2~15_combout )))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux2~15_combout ),
	.datad(\Mux2~13_combout ),
	.cin(gnd),
	.combout(\Mux2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~16 .lut_mask = 16'hBA98;
defparam \Mux2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N16
cycloneive_lcell_comb \Mux2~19 (
// Equation(s):
// \Mux2~19_combout  = (dcifimemload_24 & ((\Mux2~16_combout  & (\Mux2~18_combout )) # (!\Mux2~16_combout  & ((\Mux2~11_combout ))))) # (!dcifimemload_24 & (((\Mux2~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux2~18_combout ),
	.datac(\Mux2~11_combout ),
	.datad(\Mux2~16_combout ),
	.cin(gnd),
	.combout(\Mux2~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~19 .lut_mask = 16'hDDA0;
defparam \Mux2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N30
cycloneive_lcell_comb \regs~10 (
// Equation(s):
// \regs~10_combout  = (!\Equal0~1_combout  & \Selector3~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Equal0~1_combout ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\regs~10_combout ),
	.cout());
// synopsys translate_off
defparam \regs~10 .lut_mask = 16'h0F00;
defparam \regs~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N27
dffeas \regs[30][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][28] .is_wysiwyg = "true";
defparam \regs[30][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N1
dffeas \regs[18][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][28] .is_wysiwyg = "true";
defparam \regs[18][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N0
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[26][28]~q )) # (!dcifimemload_19 & ((\regs[18][28]~q )))))

	.dataa(\regs[26][28]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][28]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hEE30;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N26
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (dcifimemload_18 & ((\Mux35~2_combout  & ((\regs[30][28]~q ))) # (!\Mux35~2_combout  & (\regs[22][28]~q )))) # (!dcifimemload_18 & (((\Mux35~2_combout ))))

	.dataa(\regs[22][28]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[30][28]~q ),
	.datad(\Mux35~2_combout ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hF388;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N15
dffeas \regs[20][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][28] .is_wysiwyg = "true";
defparam \regs[20][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N29
dffeas \regs[28][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][28] .is_wysiwyg = "true";
defparam \regs[28][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N21
dffeas \regs[24][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][28] .is_wysiwyg = "true";
defparam \regs[24][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N19
dffeas \regs[16][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][28] .is_wysiwyg = "true";
defparam \regs[16][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N18
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[24][28]~q )) # (!dcifimemload_19 & ((\regs[16][28]~q )))))

	.dataa(dcifimemload_18),
	.datab(\regs[24][28]~q ),
	.datac(\regs[16][28]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hEE50;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N28
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (dcifimemload_18 & ((\Mux35~4_combout  & ((\regs[28][28]~q ))) # (!\Mux35~4_combout  & (\regs[20][28]~q )))) # (!dcifimemload_18 & (((\Mux35~4_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[20][28]~q ),
	.datac(\regs[28][28]~q ),
	.datad(\Mux35~4_combout ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'hF588;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N10
cycloneive_lcell_comb \Mux35~6 (
// Equation(s):
// \Mux35~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux35~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & ((\Mux35~5_combout ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux35~3_combout ),
	.datad(\Mux35~5_combout ),
	.cin(gnd),
	.combout(\Mux35~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~6 .lut_mask = 16'hB9A8;
defparam \Mux35~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N11
dffeas \regs[27][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][28] .is_wysiwyg = "true";
defparam \regs[27][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N8
cycloneive_lcell_comb \regs[31][28]~feeder (
// Equation(s):
// \regs[31][28]~feeder_combout  = \regs~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~10_combout ),
	.cin(gnd),
	.combout(\regs[31][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][28]~feeder .lut_mask = 16'hFF00;
defparam \regs[31][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N9
dffeas \regs[31][28] (
	.clk(CLK),
	.d(\regs[31][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][28] .is_wysiwyg = "true";
defparam \regs[31][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N16
cycloneive_lcell_comb \regs[19][28]~feeder (
// Equation(s):
// \regs[19][28]~feeder_combout  = \regs~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~10_combout ),
	.cin(gnd),
	.combout(\regs[19][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][28]~feeder .lut_mask = 16'hFF00;
defparam \regs[19][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N17
dffeas \regs[19][28] (
	.clk(CLK),
	.d(\regs[19][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][28] .is_wysiwyg = "true";
defparam \regs[19][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N2
cycloneive_lcell_comb \Mux35~7 (
// Equation(s):
// \Mux35~7_combout  = (dcifimemload_18 & ((\regs[23][28]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[19][28]~q  & !dcifimemload_19))))

	.dataa(\regs[23][28]~q ),
	.datab(\regs[19][28]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux35~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~7 .lut_mask = 16'hF0AC;
defparam \Mux35~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N26
cycloneive_lcell_comb \Mux35~8 (
// Equation(s):
// \Mux35~8_combout  = (dcifimemload_19 & ((\Mux35~7_combout  & ((\regs[31][28]~q ))) # (!\Mux35~7_combout  & (\regs[27][28]~q )))) # (!dcifimemload_19 & (((\Mux35~7_combout ))))

	.dataa(\regs[27][28]~q ),
	.datab(\regs[31][28]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux35~7_combout ),
	.cin(gnd),
	.combout(\Mux35~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~8 .lut_mask = 16'hCFA0;
defparam \Mux35~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N22
cycloneive_lcell_comb \regs[29][28]~feeder (
// Equation(s):
// \regs[29][28]~feeder_combout  = \regs~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[29][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[29][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N23
dffeas \regs[29][28] (
	.clk(CLK),
	.d(\regs[29][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][28] .is_wysiwyg = "true";
defparam \regs[29][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N25
dffeas \regs[25][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][28] .is_wysiwyg = "true";
defparam \regs[25][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N16
cycloneive_lcell_comb \regs[17][28]~feeder (
// Equation(s):
// \regs[17][28]~feeder_combout  = \regs~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[17][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[17][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N17
dffeas \regs[17][28] (
	.clk(CLK),
	.d(\regs[17][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][28] .is_wysiwyg = "true";
defparam \regs[17][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N18
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[21][28]~q )) # (!dcifimemload_18 & ((\regs[17][28]~q )))))

	.dataa(\regs[21][28]~q ),
	.datab(\regs[17][28]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hFA0C;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N0
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (dcifimemload_19 & ((\Mux35~0_combout  & (\regs[29][28]~q )) # (!\Mux35~0_combout  & ((\regs[25][28]~q ))))) # (!dcifimemload_19 & (((\Mux35~0_combout ))))

	.dataa(\regs[29][28]~q ),
	.datab(\regs[25][28]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux35~0_combout ),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hAFC0;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N25
dffeas \regs[14][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][28] .is_wysiwyg = "true";
defparam \regs[14][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N14
cycloneive_lcell_comb \regs[13][28]~feeder (
// Equation(s):
// \regs[13][28]~feeder_combout  = \regs~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[13][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[13][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N15
dffeas \regs[13][28] (
	.clk(CLK),
	.d(\regs[13][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][28] .is_wysiwyg = "true";
defparam \regs[13][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N5
dffeas \regs[12][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][28] .is_wysiwyg = "true";
defparam \regs[12][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N4
cycloneive_lcell_comb \Mux35~17 (
// Equation(s):
// \Mux35~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][28]~q )) # (!dcifimemload_16 & ((\regs[12][28]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[13][28]~q ),
	.datac(\regs[12][28]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux35~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~17 .lut_mask = 16'hEE50;
defparam \Mux35~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y31_N27
dffeas \regs[15][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][28] .is_wysiwyg = "true";
defparam \regs[15][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N26
cycloneive_lcell_comb \Mux35~18 (
// Equation(s):
// \Mux35~18_combout  = (\Mux35~17_combout  & (((\regs[15][28]~q ) # (!dcifimemload_17)))) # (!\Mux35~17_combout  & (\regs[14][28]~q  & ((dcifimemload_17))))

	.dataa(\regs[14][28]~q ),
	.datab(\Mux35~17_combout ),
	.datac(\regs[15][28]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux35~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~18 .lut_mask = 16'hE2CC;
defparam \Mux35~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N15
dffeas \regs[9][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][28] .is_wysiwyg = "true";
defparam \regs[9][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N3
dffeas \regs[11][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][28] .is_wysiwyg = "true";
defparam \regs[11][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N1
dffeas \regs[10][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][28] .is_wysiwyg = "true";
defparam \regs[10][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N17
dffeas \regs[8][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][28] .is_wysiwyg = "true";
defparam \regs[8][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N16
cycloneive_lcell_comb \Mux35~10 (
// Equation(s):
// \Mux35~10_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][28]~q )) # (!dcifimemload_17 & ((\regs[8][28]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][28]~q ),
	.datac(\regs[8][28]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux35~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~10 .lut_mask = 16'hEE50;
defparam \Mux35~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N2
cycloneive_lcell_comb \Mux35~11 (
// Equation(s):
// \Mux35~11_combout  = (dcifimemload_16 & ((\Mux35~10_combout  & ((\regs[11][28]~q ))) # (!\Mux35~10_combout  & (\regs[9][28]~q )))) # (!dcifimemload_16 & (((\Mux35~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][28]~q ),
	.datac(\regs[11][28]~q ),
	.datad(\Mux35~10_combout ),
	.cin(gnd),
	.combout(\Mux35~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~11 .lut_mask = 16'hF588;
defparam \Mux35~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y32_N19
dffeas \regs[2][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][28] .is_wysiwyg = "true";
defparam \regs[2][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N1
dffeas \regs[1][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][28] .is_wysiwyg = "true";
defparam \regs[1][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N0
cycloneive_lcell_comb \Mux35~14 (
// Equation(s):
// \Mux35~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][28]~q )) # (!dcifimemload_17 & ((\regs[1][28]~q )))))

	.dataa(\regs[3][28]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][28]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux35~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~14 .lut_mask = 16'h88C0;
defparam \Mux35~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N18
cycloneive_lcell_comb \Mux35~15 (
// Equation(s):
// \Mux35~15_combout  = (\Mux35~14_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][28]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[2][28]~q ),
	.datad(\Mux35~14_combout ),
	.cin(gnd),
	.combout(\Mux35~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~15 .lut_mask = 16'hFF20;
defparam \Mux35~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N13
dffeas \regs[6][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][28] .is_wysiwyg = "true";
defparam \regs[6][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N15
dffeas \regs[7][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][28] .is_wysiwyg = "true";
defparam \regs[7][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N13
dffeas \regs[4][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][28] .is_wysiwyg = "true";
defparam \regs[4][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N12
cycloneive_lcell_comb \Mux35~12 (
// Equation(s):
// \Mux35~12_combout  = (dcifimemload_16 & ((\regs[5][28]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][28]~q  & !dcifimemload_17))))

	.dataa(\regs[5][28]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][28]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux35~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~12 .lut_mask = 16'hCCB8;
defparam \Mux35~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N14
cycloneive_lcell_comb \Mux35~13 (
// Equation(s):
// \Mux35~13_combout  = (dcifimemload_17 & ((\Mux35~12_combout  & ((\regs[7][28]~q ))) # (!\Mux35~12_combout  & (\regs[6][28]~q )))) # (!dcifimemload_17 & (((\Mux35~12_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][28]~q ),
	.datac(\regs[7][28]~q ),
	.datad(\Mux35~12_combout ),
	.cin(gnd),
	.combout(\Mux35~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~13 .lut_mask = 16'hF588;
defparam \Mux35~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N16
cycloneive_lcell_comb \Mux35~16 (
// Equation(s):
// \Mux35~16_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux35~13_combout ))) # (!dcifimemload_18 & (\Mux35~15_combout ))))

	.dataa(\Mux35~15_combout ),
	.datab(dcifimemload_19),
	.datac(dcifimemload_18),
	.datad(\Mux35~13_combout ),
	.cin(gnd),
	.combout(\Mux35~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~16 .lut_mask = 16'hF2C2;
defparam \Mux35~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N20
cycloneive_lcell_comb \Mux3~17 (
// Equation(s):
// \Mux3~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\regs[13][28]~q ))) # (!dcifimemload_21 & (\regs[12][28]~q ))))

	.dataa(\regs[12][28]~q ),
	.datab(\regs[13][28]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux3~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~17 .lut_mask = 16'hFC0A;
defparam \Mux3~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N24
cycloneive_lcell_comb \Mux3~18 (
// Equation(s):
// \Mux3~18_combout  = (dcifimemload_22 & ((\Mux3~17_combout  & (\regs[15][28]~q )) # (!\Mux3~17_combout  & ((\regs[14][28]~q ))))) # (!dcifimemload_22 & (((\Mux3~17_combout ))))

	.dataa(\regs[15][28]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[14][28]~q ),
	.datad(\Mux3~17_combout ),
	.cin(gnd),
	.combout(\Mux3~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~18 .lut_mask = 16'hBBC0;
defparam \Mux3~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \Mux3~12 (
// Equation(s):
// \Mux3~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][28]~q ))) # (!dcifimemload_22 & (\regs[8][28]~q ))))

	.dataa(\regs[8][28]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[10][28]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux3~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~12 .lut_mask = 16'hFC22;
defparam \Mux3~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N24
cycloneive_lcell_comb \Mux3~13 (
// Equation(s):
// \Mux3~13_combout  = (dcifimemload_21 & ((\Mux3~12_combout  & (\regs[11][28]~q )) # (!\Mux3~12_combout  & ((\regs[9][28]~q ))))) # (!dcifimemload_21 & (((\Mux3~12_combout ))))

	.dataa(\regs[11][28]~q ),
	.datab(\regs[9][28]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux3~12_combout ),
	.cin(gnd),
	.combout(\Mux3~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~13 .lut_mask = 16'hAFC0;
defparam \Mux3~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N0
cycloneive_lcell_comb \regs[3][28]~feeder (
// Equation(s):
// \regs[3][28]~feeder_combout  = \regs~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~10_combout ),
	.cin(gnd),
	.combout(\regs[3][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][28]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N1
dffeas \regs[3][28] (
	.clk(CLK),
	.d(\regs[3][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][28] .is_wysiwyg = "true";
defparam \regs[3][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N18
cycloneive_lcell_comb \Mux3~14 (
// Equation(s):
// \Mux3~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][28]~q ))) # (!dcifimemload_22 & (\regs[1][28]~q ))))

	.dataa(\regs[1][28]~q ),
	.datab(\regs[3][28]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux3~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~14 .lut_mask = 16'hC0A0;
defparam \Mux3~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N16
cycloneive_lcell_comb \Mux3~15 (
// Equation(s):
// \Mux3~15_combout  = (\Mux3~14_combout ) # ((\regs[2][28]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\regs[2][28]~q ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux3~14_combout ),
	.cin(gnd),
	.combout(\Mux3~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~15 .lut_mask = 16'hFF08;
defparam \Mux3~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N26
cycloneive_lcell_comb \Mux3~16 (
// Equation(s):
// \Mux3~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & (\Mux3~13_combout )) # (!dcifimemload_24 & ((\Mux3~15_combout )))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux3~13_combout ),
	.datad(\Mux3~15_combout ),
	.cin(gnd),
	.combout(\Mux3~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~16 .lut_mask = 16'hD9C8;
defparam \Mux3~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N7
dffeas \regs[5][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][28] .is_wysiwyg = "true";
defparam \regs[5][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N6
cycloneive_lcell_comb \Mux3~10 (
// Equation(s):
// \Mux3~10_combout  = (dcifimemload_21 & (((\regs[5][28]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][28]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][28]~q ),
	.datac(\regs[5][28]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~10 .lut_mask = 16'hAAE4;
defparam \Mux3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N12
cycloneive_lcell_comb \Mux3~11 (
// Equation(s):
// \Mux3~11_combout  = (dcifimemload_22 & ((\Mux3~10_combout  & (\regs[7][28]~q )) # (!\Mux3~10_combout  & ((\regs[6][28]~q ))))) # (!dcifimemload_22 & (((\Mux3~10_combout ))))

	.dataa(\regs[7][28]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[6][28]~q ),
	.datad(\Mux3~10_combout ),
	.cin(gnd),
	.combout(\Mux3~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~11 .lut_mask = 16'hBBC0;
defparam \Mux3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N4
cycloneive_lcell_comb \Mux3~19 (
// Equation(s):
// \Mux3~19_combout  = (dcifimemload_23 & ((\Mux3~16_combout  & (\Mux3~18_combout )) # (!\Mux3~16_combout  & ((\Mux3~11_combout ))))) # (!dcifimemload_23 & (((\Mux3~16_combout ))))

	.dataa(\Mux3~18_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux3~16_combout ),
	.datad(\Mux3~11_combout ),
	.cin(gnd),
	.combout(\Mux3~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~19 .lut_mask = 16'hBCB0;
defparam \Mux3~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N30
cycloneive_lcell_comb \regs[23][28]~feeder (
// Equation(s):
// \regs[23][28]~feeder_combout  = \regs~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~10_combout ),
	.cin(gnd),
	.combout(\regs[23][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][28]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N31
dffeas \regs[23][28] (
	.clk(CLK),
	.d(\regs[23][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][28] .is_wysiwyg = "true";
defparam \regs[23][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N10
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (dcifimemload_24 & (((\regs[27][28]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[19][28]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[19][28]~q ),
	.datac(\regs[27][28]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hAAE4;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N4
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (dcifimemload_23 & ((\Mux3~7_combout  & (\regs[31][28]~q )) # (!\Mux3~7_combout  & ((\regs[23][28]~q ))))) # (!dcifimemload_23 & (((\Mux3~7_combout ))))

	.dataa(\regs[31][28]~q ),
	.datab(\regs[23][28]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux3~7_combout ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hAFC0;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N30
cycloneive_lcell_comb \regs[21][28]~feeder (
// Equation(s):
// \regs[21][28]~feeder_combout  = \regs~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[21][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[21][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y31_N31
dffeas \regs[21][28] (
	.clk(CLK),
	.d(\regs[21][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][28] .is_wysiwyg = "true";
defparam \regs[21][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N24
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (dcifimemload_24 & (((\regs[25][28]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[17][28]~q  & ((!dcifimemload_23))))

	.dataa(\regs[17][28]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[25][28]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hCCE2;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N20
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (dcifimemload_23 & ((\Mux3~0_combout  & (\regs[29][28]~q )) # (!\Mux3~0_combout  & ((\regs[21][28]~q ))))) # (!dcifimemload_23 & (((\Mux3~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[29][28]~q ),
	.datac(\regs[21][28]~q ),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hDDA0;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N14
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[20][28]~q ))) # (!dcifimemload_23 & (\regs[16][28]~q ))))

	.dataa(dcifimemload_24),
	.datab(\regs[16][28]~q ),
	.datac(\regs[20][28]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hFA44;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N20
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (dcifimemload_24 & ((\Mux3~4_combout  & (\regs[28][28]~q )) # (!\Mux3~4_combout  & ((\regs[24][28]~q ))))) # (!dcifimemload_24 & (((\Mux3~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[28][28]~q ),
	.datac(\regs[24][28]~q ),
	.datad(\Mux3~4_combout ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hDDA0;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N22
cycloneive_lcell_comb \regs[26][28]~feeder (
// Equation(s):
// \regs[26][28]~feeder_combout  = \regs~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[26][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[26][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N23
dffeas \regs[26][28] (
	.clk(CLK),
	.d(\regs[26][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][28] .is_wysiwyg = "true";
defparam \regs[26][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N1
dffeas \regs[22][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][28] .is_wysiwyg = "true";
defparam \regs[22][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N0
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (dcifimemload_23 & (((\regs[22][28]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[18][28]~q  & ((!dcifimemload_24))))

	.dataa(\regs[18][28]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[22][28]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hCCE2;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N8
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (dcifimemload_24 & ((\Mux3~2_combout  & (\regs[30][28]~q )) # (!\Mux3~2_combout  & ((\regs[26][28]~q ))))) # (!dcifimemload_24 & (((\Mux3~2_combout ))))

	.dataa(\regs[30][28]~q ),
	.datab(\regs[26][28]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux3~2_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hAFC0;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N12
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux3~3_combout ))) # (!dcifimemload_22 & (\Mux3~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux3~5_combout ),
	.datad(\Mux3~3_combout ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hDC98;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N2
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// \Mux3~9_combout  = (dcifimemload_21 & ((\Mux3~6_combout  & (\Mux3~8_combout )) # (!\Mux3~6_combout  & ((\Mux3~1_combout ))))) # (!dcifimemload_21 & (((\Mux3~6_combout ))))

	.dataa(\Mux3~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux3~1_combout ),
	.datad(\Mux3~6_combout ),
	.cin(gnd),
	.combout(\Mux3~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hBBC0;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N8
cycloneive_lcell_comb \regs~11 (
// Equation(s):
// \regs~11_combout  = (cuifRegSel_11 & ((dcifimemload_11) # ((!cuifRegSel_0)))) # (!cuifRegSel_11 & (((cuifRegSel_0 & ramiframload_271))))

	.dataa(cuifRegSel_11),
	.datab(dcifimemload_11),
	.datac(cuifRegSel_0),
	.datad(ramiframload_27),
	.cin(gnd),
	.combout(\regs~11_combout ),
	.cout());
// synopsys translate_off
defparam \regs~11 .lut_mask = 16'hDA8A;
defparam \regs~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N22
cycloneive_lcell_comb \regs~13 (
// Equation(s):
// \regs~13_combout  = (!\Equal0~1_combout  & ((\regs~12_combout  & ((\regs~11_combout ))) # (!\regs~12_combout  & (Mux410 & !\regs~11_combout ))))

	.dataa(\regs~12_combout ),
	.datab(\Equal0~1_combout ),
	.datac(Mux410),
	.datad(\regs~11_combout ),
	.cin(gnd),
	.combout(\regs~13_combout ),
	.cout());
// synopsys translate_off
defparam \regs~13 .lut_mask = 16'h2210;
defparam \regs~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N10
cycloneive_lcell_comb \regs[20][27]~feeder (
// Equation(s):
// \regs[20][27]~feeder_combout  = \regs~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[20][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[20][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N11
dffeas \regs[20][27] (
	.clk(CLK),
	.d(\regs[20][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][27] .is_wysiwyg = "true";
defparam \regs[20][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N3
dffeas \regs[16][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][27] .is_wysiwyg = "true";
defparam \regs[16][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N2
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (dcifimemload_18 & ((\regs[20][27]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[16][27]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[20][27]~q ),
	.datac(\regs[16][27]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'hAAD8;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N5
dffeas \regs[28][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][27] .is_wysiwyg = "true";
defparam \regs[28][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N4
cycloneive_lcell_comb \Mux36~5 (
// Equation(s):
// \Mux36~5_combout  = (\Mux36~4_combout  & (((\regs[28][27]~q ) # (!dcifimemload_19)))) # (!\Mux36~4_combout  & (\regs[24][27]~q  & ((dcifimemload_19))))

	.dataa(\regs[24][27]~q ),
	.datab(\Mux36~4_combout ),
	.datac(\regs[28][27]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux36~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~5 .lut_mask = 16'hE2CC;
defparam \Mux36~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N13
dffeas \regs[30][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][27] .is_wysiwyg = "true";
defparam \regs[30][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N11
dffeas \regs[18][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][27] .is_wysiwyg = "true";
defparam \regs[18][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N10
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (dcifimemload_18 & ((\regs[22][27]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[18][27]~q  & !dcifimemload_19))))

	.dataa(\regs[22][27]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][27]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'hCCB8;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N12
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (dcifimemload_19 & ((\Mux36~2_combout  & ((\regs[30][27]~q ))) # (!\Mux36~2_combout  & (\regs[26][27]~q )))) # (!dcifimemload_19 & (((\Mux36~2_combout ))))

	.dataa(\regs[26][27]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[30][27]~q ),
	.datad(\Mux36~2_combout ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hF388;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N6
cycloneive_lcell_comb \Mux36~6 (
// Equation(s):
// \Mux36~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux36~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux36~5_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux36~5_combout ),
	.datad(\Mux36~3_combout ),
	.cin(gnd),
	.combout(\Mux36~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~6 .lut_mask = 16'hBA98;
defparam \Mux36~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N12
cycloneive_lcell_comb \regs[23][27]~feeder (
// Equation(s):
// \regs[23][27]~feeder_combout  = \regs~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~13_combout ),
	.cin(gnd),
	.combout(\regs[23][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][27]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N13
dffeas \regs[23][27] (
	.clk(CLK),
	.d(\regs[23][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][27] .is_wysiwyg = "true";
defparam \regs[23][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N20
cycloneive_lcell_comb \regs[31][27]~feeder (
// Equation(s):
// \regs[31][27]~feeder_combout  = \regs~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[31][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[31][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N21
dffeas \regs[31][27] (
	.clk(CLK),
	.d(\regs[31][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][27] .is_wysiwyg = "true";
defparam \regs[31][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N31
dffeas \regs[27][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][27] .is_wysiwyg = "true";
defparam \regs[27][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N10
cycloneive_lcell_comb \Mux36~7 (
// Equation(s):
// \Mux36~7_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[27][27]~q ))) # (!dcifimemload_19 & (\regs[19][27]~q ))))

	.dataa(\regs[19][27]~q ),
	.datab(\regs[27][27]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux36~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~7 .lut_mask = 16'hFC0A;
defparam \Mux36~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N14
cycloneive_lcell_comb \Mux36~8 (
// Equation(s):
// \Mux36~8_combout  = (dcifimemload_18 & ((\Mux36~7_combout  & ((\regs[31][27]~q ))) # (!\Mux36~7_combout  & (\regs[23][27]~q )))) # (!dcifimemload_18 & (((\Mux36~7_combout ))))

	.dataa(\regs[23][27]~q ),
	.datab(\regs[31][27]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux36~7_combout ),
	.cin(gnd),
	.combout(\Mux36~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~8 .lut_mask = 16'hCFA0;
defparam \Mux36~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N20
cycloneive_lcell_comb \regs[21][27]~feeder (
// Equation(s):
// \regs[21][27]~feeder_combout  = \regs~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[21][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[21][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N21
dffeas \regs[21][27] (
	.clk(CLK),
	.d(\regs[21][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][27] .is_wysiwyg = "true";
defparam \regs[21][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N29
dffeas \regs[29][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][27] .is_wysiwyg = "true";
defparam \regs[29][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N17
dffeas \regs[25][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][27] .is_wysiwyg = "true";
defparam \regs[25][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N31
dffeas \regs[17][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][27] .is_wysiwyg = "true";
defparam \regs[17][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N30
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[25][27]~q )) # (!dcifimemload_19 & ((\regs[17][27]~q )))))

	.dataa(dcifimemload_18),
	.datab(\regs[25][27]~q ),
	.datac(\regs[17][27]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hEE50;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N28
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (dcifimemload_18 & ((\Mux36~0_combout  & ((\regs[29][27]~q ))) # (!\Mux36~0_combout  & (\regs[21][27]~q )))) # (!dcifimemload_18 & (((\Mux36~0_combout ))))

	.dataa(\regs[21][27]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[29][27]~q ),
	.datad(\Mux36~0_combout ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hF388;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N17
dffeas \regs[6][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][27] .is_wysiwyg = "true";
defparam \regs[6][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N23
dffeas \regs[7][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][27] .is_wysiwyg = "true";
defparam \regs[7][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N17
dffeas \regs[4][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][27] .is_wysiwyg = "true";
defparam \regs[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N16
cycloneive_lcell_comb \Mux36~10 (
// Equation(s):
// \Mux36~10_combout  = (dcifimemload_16 & ((\regs[5][27]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][27]~q  & !dcifimemload_17))))

	.dataa(\regs[5][27]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][27]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux36~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~10 .lut_mask = 16'hCCB8;
defparam \Mux36~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N22
cycloneive_lcell_comb \Mux36~11 (
// Equation(s):
// \Mux36~11_combout  = (dcifimemload_17 & ((\Mux36~10_combout  & ((\regs[7][27]~q ))) # (!\Mux36~10_combout  & (\regs[6][27]~q )))) # (!dcifimemload_17 & (((\Mux36~10_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][27]~q ),
	.datac(\regs[7][27]~q ),
	.datad(\Mux36~10_combout ),
	.cin(gnd),
	.combout(\Mux36~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~11 .lut_mask = 16'hF588;
defparam \Mux36~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N7
dffeas \regs[2][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][27] .is_wysiwyg = "true";
defparam \regs[2][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N29
dffeas \regs[3][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][27] .is_wysiwyg = "true";
defparam \regs[3][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N25
dffeas \regs[1][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][27] .is_wysiwyg = "true";
defparam \regs[1][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N24
cycloneive_lcell_comb \Mux36~14 (
// Equation(s):
// \Mux36~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][27]~q )) # (!dcifimemload_17 & ((\regs[1][27]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[3][27]~q ),
	.datac(\regs[1][27]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux36~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~14 .lut_mask = 16'h88A0;
defparam \Mux36~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N6
cycloneive_lcell_comb \Mux36~15 (
// Equation(s):
// \Mux36~15_combout  = (\Mux36~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][27]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][27]~q ),
	.datad(\Mux36~14_combout ),
	.cin(gnd),
	.combout(\Mux36~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~15 .lut_mask = 16'hFF40;
defparam \Mux36~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N9
dffeas \regs[8][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][27] .is_wysiwyg = "true";
defparam \regs[8][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \regs[10][27]~feeder (
// Equation(s):
// \regs[10][27]~feeder_combout  = \regs~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~13_combout ),
	.cin(gnd),
	.combout(\regs[10][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[10][27]~feeder .lut_mask = 16'hFF00;
defparam \regs[10][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N11
dffeas \regs[10][27] (
	.clk(CLK),
	.d(\regs[10][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][27] .is_wysiwyg = "true";
defparam \regs[10][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N8
cycloneive_lcell_comb \Mux36~12 (
// Equation(s):
// \Mux36~12_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\regs[10][27]~q )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\regs[8][27]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[8][27]~q ),
	.datad(\regs[10][27]~q ),
	.cin(gnd),
	.combout(\Mux36~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~12 .lut_mask = 16'hBA98;
defparam \Mux36~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N27
dffeas \regs[11][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][27] .is_wysiwyg = "true";
defparam \regs[11][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N3
dffeas \regs[9][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][27] .is_wysiwyg = "true";
defparam \regs[9][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N26
cycloneive_lcell_comb \Mux36~13 (
// Equation(s):
// \Mux36~13_combout  = (dcifimemload_16 & ((\Mux36~12_combout  & (\regs[11][27]~q )) # (!\Mux36~12_combout  & ((\regs[9][27]~q ))))) # (!dcifimemload_16 & (\Mux36~12_combout ))

	.dataa(dcifimemload_16),
	.datab(\Mux36~12_combout ),
	.datac(\regs[11][27]~q ),
	.datad(\regs[9][27]~q ),
	.cin(gnd),
	.combout(\Mux36~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~13 .lut_mask = 16'hE6C4;
defparam \Mux36~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N30
cycloneive_lcell_comb \Mux36~16 (
// Equation(s):
// \Mux36~16_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & ((\Mux36~13_combout ))) # (!dcifimemload_19 & (\Mux36~15_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux36~15_combout ),
	.datad(\Mux36~13_combout ),
	.cin(gnd),
	.combout(\Mux36~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~16 .lut_mask = 16'hDC98;
defparam \Mux36~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N11
dffeas \regs[14][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][27] .is_wysiwyg = "true";
defparam \regs[14][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N11
dffeas \regs[15][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][27] .is_wysiwyg = "true";
defparam \regs[15][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N1
dffeas \regs[13][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][27] .is_wysiwyg = "true";
defparam \regs[13][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N17
dffeas \regs[12][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][27] .is_wysiwyg = "true";
defparam \regs[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N16
cycloneive_lcell_comb \Mux36~17 (
// Equation(s):
// \Mux36~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][27]~q )) # (!dcifimemload_16 & ((\regs[12][27]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[13][27]~q ),
	.datac(\regs[12][27]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux36~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~17 .lut_mask = 16'hEE50;
defparam \Mux36~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N10
cycloneive_lcell_comb \Mux36~18 (
// Equation(s):
// \Mux36~18_combout  = (dcifimemload_17 & ((\Mux36~17_combout  & ((\regs[15][27]~q ))) # (!\Mux36~17_combout  & (\regs[14][27]~q )))) # (!dcifimemload_17 & (((\Mux36~17_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[14][27]~q ),
	.datac(\regs[15][27]~q ),
	.datad(\Mux36~17_combout ),
	.cin(gnd),
	.combout(\Mux36~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~18 .lut_mask = 16'hF588;
defparam \Mux36~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N12
cycloneive_lcell_comb \regs[19][27]~feeder (
// Equation(s):
// \regs[19][27]~feeder_combout  = \regs~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[19][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[19][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N13
dffeas \regs[19][27] (
	.clk(CLK),
	.d(\regs[19][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][27] .is_wysiwyg = "true";
defparam \regs[19][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N22
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[23][27]~q )) # (!dcifimemload_23 & ((\regs[19][27]~q )))))

	.dataa(\regs[23][27]~q ),
	.datab(\regs[19][27]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hFA0C;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N30
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (dcifimemload_24 & ((\Mux4~7_combout  & (\regs[31][27]~q )) # (!\Mux4~7_combout  & ((\regs[27][27]~q ))))) # (!dcifimemload_24 & (((\Mux4~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[31][27]~q ),
	.datac(\regs[27][27]~q ),
	.datad(\Mux4~7_combout ),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'hDDA0;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N12
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[21][27]~q ))) # (!dcifimemload_23 & (\regs[17][27]~q ))))

	.dataa(\regs[17][27]~q ),
	.datab(\regs[21][27]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hFC0A;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N16
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (dcifimemload_24 & ((\Mux4~0_combout  & (\regs[29][27]~q )) # (!\Mux4~0_combout  & ((\regs[25][27]~q ))))) # (!dcifimemload_24 & (((\Mux4~0_combout ))))

	.dataa(\regs[29][27]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[25][27]~q ),
	.datad(\Mux4~0_combout ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hBBC0;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N0
cycloneive_lcell_comb \regs[22][27]~feeder (
// Equation(s):
// \regs[22][27]~feeder_combout  = \regs~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[22][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[22][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N1
dffeas \regs[22][27] (
	.clk(CLK),
	.d(\regs[22][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][27] .is_wysiwyg = "true";
defparam \regs[22][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N7
dffeas \regs[26][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][27] .is_wysiwyg = "true";
defparam \regs[26][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N6
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\regs[26][27]~q ))) # (!dcifimemload_24 & (\regs[18][27]~q ))))

	.dataa(dcifimemload_23),
	.datab(\regs[18][27]~q ),
	.datac(\regs[26][27]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hFA44;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N12
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (dcifimemload_23 & ((\Mux4~2_combout  & (\regs[30][27]~q )) # (!\Mux4~2_combout  & ((\regs[22][27]~q ))))) # (!dcifimemload_23 & (((\Mux4~2_combout ))))

	.dataa(\regs[30][27]~q ),
	.datab(\regs[22][27]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux4~2_combout ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hAFC0;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N19
dffeas \regs[24][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][27] .is_wysiwyg = "true";
defparam \regs[24][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N18
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (dcifimemload_24 & (((\regs[24][27]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[16][27]~q  & ((!dcifimemload_23))))

	.dataa(\regs[16][27]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[24][27]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hCCE2;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N22
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (dcifimemload_23 & ((\Mux4~4_combout  & ((\regs[28][27]~q ))) # (!\Mux4~4_combout  & (\regs[20][27]~q )))) # (!dcifimemload_23 & (((\Mux4~4_combout ))))

	.dataa(\regs[20][27]~q ),
	.datab(\regs[28][27]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux4~4_combout ),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hCFA0;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N12
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux4~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux4~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux4~3_combout ),
	.datad(\Mux4~5_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hB9A8;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N30
cycloneive_lcell_comb \Mux4~9 (
// Equation(s):
// \Mux4~9_combout  = (dcifimemload_21 & ((\Mux4~6_combout  & (\Mux4~8_combout )) # (!\Mux4~6_combout  & ((\Mux4~1_combout ))))) # (!dcifimemload_21 & (((\Mux4~6_combout ))))

	.dataa(\Mux4~8_combout ),
	.datab(\Mux4~1_combout ),
	.datac(dcifimemload_21),
	.datad(\Mux4~6_combout ),
	.cin(gnd),
	.combout(\Mux4~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~9 .lut_mask = 16'hAFC0;
defparam \Mux4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N0
cycloneive_lcell_comb \Mux4~17 (
// Equation(s):
// \Mux4~17_combout  = (dcifimemload_21 & (((\regs[13][27]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][27]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][27]~q ),
	.datac(\regs[13][27]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux4~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~17 .lut_mask = 16'hAAE4;
defparam \Mux4~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N10
cycloneive_lcell_comb \Mux4~18 (
// Equation(s):
// \Mux4~18_combout  = (dcifimemload_22 & ((\Mux4~17_combout  & (\regs[15][27]~q )) # (!\Mux4~17_combout  & ((\regs[14][27]~q ))))) # (!dcifimemload_22 & (((\Mux4~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][27]~q ),
	.datac(\regs[14][27]~q ),
	.datad(\Mux4~17_combout ),
	.cin(gnd),
	.combout(\Mux4~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~18 .lut_mask = 16'hDDA0;
defparam \Mux4~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N24
cycloneive_lcell_comb \Mux4~10 (
// Equation(s):
// \Mux4~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\regs[10][27]~q )) # (!dcifimemload_22 & ((\regs[8][27]~q )))))

	.dataa(\regs[10][27]~q ),
	.datab(\regs[8][27]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~10 .lut_mask = 16'hFA0C;
defparam \Mux4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N2
cycloneive_lcell_comb \Mux4~11 (
// Equation(s):
// \Mux4~11_combout  = (dcifimemload_21 & ((\Mux4~10_combout  & (\regs[11][27]~q )) # (!\Mux4~10_combout  & ((\regs[9][27]~q ))))) # (!dcifimemload_21 & (((\Mux4~10_combout ))))

	.dataa(\regs[11][27]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[9][27]~q ),
	.datad(\Mux4~10_combout ),
	.cin(gnd),
	.combout(\Mux4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~11 .lut_mask = 16'hBBC0;
defparam \Mux4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N28
cycloneive_lcell_comb \Mux4~14 (
// Equation(s):
// \Mux4~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][27]~q ))) # (!dcifimemload_22 & (\regs[1][27]~q ))))

	.dataa(\regs[1][27]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[3][27]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux4~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~14 .lut_mask = 16'hC088;
defparam \Mux4~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N8
cycloneive_lcell_comb \Mux4~15 (
// Equation(s):
// \Mux4~15_combout  = (\Mux4~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][27]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[2][27]~q ),
	.datad(\Mux4~14_combout ),
	.cin(gnd),
	.combout(\Mux4~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~15 .lut_mask = 16'hFF20;
defparam \Mux4~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N19
dffeas \regs[5][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][27] .is_wysiwyg = "true";
defparam \regs[5][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N18
cycloneive_lcell_comb \Mux4~12 (
// Equation(s):
// \Mux4~12_combout  = (dcifimemload_21 & (((\regs[5][27]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][27]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][27]~q ),
	.datac(\regs[5][27]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux4~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~12 .lut_mask = 16'hAAE4;
defparam \Mux4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N16
cycloneive_lcell_comb \Mux4~13 (
// Equation(s):
// \Mux4~13_combout  = (dcifimemload_22 & ((\Mux4~12_combout  & (\regs[7][27]~q )) # (!\Mux4~12_combout  & ((\regs[6][27]~q ))))) # (!dcifimemload_22 & (((\Mux4~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[7][27]~q ),
	.datac(\regs[6][27]~q ),
	.datad(\Mux4~12_combout ),
	.cin(gnd),
	.combout(\Mux4~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~13 .lut_mask = 16'hDDA0;
defparam \Mux4~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N18
cycloneive_lcell_comb \Mux4~16 (
// Equation(s):
// \Mux4~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux4~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & (\Mux4~15_combout )))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux4~15_combout ),
	.datad(\Mux4~13_combout ),
	.cin(gnd),
	.combout(\Mux4~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~16 .lut_mask = 16'hBA98;
defparam \Mux4~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N24
cycloneive_lcell_comb \Mux4~19 (
// Equation(s):
// \Mux4~19_combout  = (dcifimemload_24 & ((\Mux4~16_combout  & (\Mux4~18_combout )) # (!\Mux4~16_combout  & ((\Mux4~11_combout ))))) # (!dcifimemload_24 & (((\Mux4~16_combout ))))

	.dataa(\Mux4~18_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux4~11_combout ),
	.datad(\Mux4~16_combout ),
	.cin(gnd),
	.combout(\Mux4~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~19 .lut_mask = 16'hBBC0;
defparam \Mux4~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N24
cycloneive_lcell_comb \regs~14 (
// Equation(s):
// \regs~14_combout  = (cuifRegSel_11 & ((cuifRegSel_0 & (dcifimemload_10)) # (!cuifRegSel_0 & ((\Add1~48_combout ))))) # (!cuifRegSel_11 & (cuifRegSel_0))

	.dataa(cuifRegSel_11),
	.datab(cuifRegSel_0),
	.datac(dcifimemload_10),
	.datad(Add116),
	.cin(gnd),
	.combout(\regs~14_combout ),
	.cout());
// synopsys translate_off
defparam \regs~14 .lut_mask = 16'hE6C4;
defparam \regs~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N12
cycloneive_lcell_comb \regs~16 (
// Equation(s):
// \regs~16_combout  = (!\Equal0~1_combout  & ((\regs~15_combout  & ((\regs~14_combout ))) # (!\regs~15_combout  & (Mux510 & !\regs~14_combout ))))

	.dataa(\regs~15_combout ),
	.datab(Mux510),
	.datac(\regs~14_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\regs~16_combout ),
	.cout());
// synopsys translate_off
defparam \regs~16 .lut_mask = 16'h00A4;
defparam \regs~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N19
dffeas \regs[20][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][26] .is_wysiwyg = "true";
defparam \regs[20][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N15
dffeas \regs[28][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][26] .is_wysiwyg = "true";
defparam \regs[28][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N1
dffeas \regs[24][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][26] .is_wysiwyg = "true";
defparam \regs[24][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N29
dffeas \regs[16][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][26] .is_wysiwyg = "true";
defparam \regs[16][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N28
cycloneive_lcell_comb \Mux37~4 (
// Equation(s):
// \Mux37~4_combout  = (dcifimemload_19 & ((\regs[24][26]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\regs[16][26]~q  & !dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\regs[24][26]~q ),
	.datac(\regs[16][26]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux37~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~4 .lut_mask = 16'hAAD8;
defparam \Mux37~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N14
cycloneive_lcell_comb \Mux37~5 (
// Equation(s):
// \Mux37~5_combout  = (dcifimemload_18 & ((\Mux37~4_combout  & ((\regs[28][26]~q ))) # (!\Mux37~4_combout  & (\regs[20][26]~q )))) # (!dcifimemload_18 & (((\Mux37~4_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[20][26]~q ),
	.datac(\regs[28][26]~q ),
	.datad(\Mux37~4_combout ),
	.cin(gnd),
	.combout(\Mux37~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~5 .lut_mask = 16'hF588;
defparam \Mux37~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N21
dffeas \regs[30][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][26] .is_wysiwyg = "true";
defparam \regs[30][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N7
dffeas \regs[22][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][26] .is_wysiwyg = "true";
defparam \regs[22][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N20
cycloneive_lcell_comb \Mux37~3 (
// Equation(s):
// \Mux37~3_combout  = (\Mux37~2_combout  & (((\regs[30][26]~q )) # (!dcifimemload_18))) # (!\Mux37~2_combout  & (dcifimemload_18 & ((\regs[22][26]~q ))))

	.dataa(\Mux37~2_combout ),
	.datab(dcifimemload_18),
	.datac(\regs[30][26]~q ),
	.datad(\regs[22][26]~q ),
	.cin(gnd),
	.combout(\Mux37~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~3 .lut_mask = 16'hE6A2;
defparam \Mux37~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N20
cycloneive_lcell_comb \Mux37~6 (
// Equation(s):
// \Mux37~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux37~3_combout ))) # (!dcifimemload_17 & (\Mux37~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux37~5_combout ),
	.datad(\Mux37~3_combout ),
	.cin(gnd),
	.combout(\Mux37~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~6 .lut_mask = 16'hDC98;
defparam \Mux37~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N20
cycloneive_lcell_comb \regs[27][26]~feeder (
// Equation(s):
// \regs[27][26]~feeder_combout  = \regs~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~16_combout ),
	.cin(gnd),
	.combout(\regs[27][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][26]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N21
dffeas \regs[27][26] (
	.clk(CLK),
	.d(\regs[27][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][26] .is_wysiwyg = "true";
defparam \regs[27][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N1
dffeas \regs[31][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][26] .is_wysiwyg = "true";
defparam \regs[31][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N17
dffeas \regs[23][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][26] .is_wysiwyg = "true";
defparam \regs[23][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N7
dffeas \regs[19][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][26] .is_wysiwyg = "true";
defparam \regs[19][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N6
cycloneive_lcell_comb \Mux37~7 (
// Equation(s):
// \Mux37~7_combout  = (dcifimemload_18 & ((\regs[23][26]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[19][26]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[23][26]~q ),
	.datac(\regs[19][26]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux37~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~7 .lut_mask = 16'hAAD8;
defparam \Mux37~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N0
cycloneive_lcell_comb \Mux37~8 (
// Equation(s):
// \Mux37~8_combout  = (dcifimemload_19 & ((\Mux37~7_combout  & ((\regs[31][26]~q ))) # (!\Mux37~7_combout  & (\regs[27][26]~q )))) # (!dcifimemload_19 & (((\Mux37~7_combout ))))

	.dataa(\regs[27][26]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[31][26]~q ),
	.datad(\Mux37~7_combout ),
	.cin(gnd),
	.combout(\Mux37~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~8 .lut_mask = 16'hF388;
defparam \Mux37~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N13
dffeas \regs[25][26] (
	.clk(CLK),
	.d(\regs~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][26] .is_wysiwyg = "true";
defparam \regs[25][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N15
dffeas \regs[29][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][26] .is_wysiwyg = "true";
defparam \regs[29][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N26
cycloneive_lcell_comb \regs[21][26]~feeder (
// Equation(s):
// \regs[21][26]~feeder_combout  = \regs~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~16_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[21][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][26]~feeder .lut_mask = 16'hF0F0;
defparam \regs[21][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N27
dffeas \regs[21][26] (
	.clk(CLK),
	.d(\regs[21][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][26] .is_wysiwyg = "true";
defparam \regs[21][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N5
dffeas \regs[17][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][26] .is_wysiwyg = "true";
defparam \regs[17][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N4
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[21][26]~q )) # (!dcifimemload_18 & ((\regs[17][26]~q )))))

	.dataa(dcifimemload_19),
	.datab(\regs[21][26]~q ),
	.datac(\regs[17][26]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hEE50;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N14
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (dcifimemload_19 & ((\Mux37~0_combout  & ((\regs[29][26]~q ))) # (!\Mux37~0_combout  & (\regs[25][26]~q )))) # (!dcifimemload_19 & (((\Mux37~0_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[25][26]~q ),
	.datac(\regs[29][26]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hF588;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N9
dffeas \regs[9][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][26] .is_wysiwyg = "true";
defparam \regs[9][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N31
dffeas \regs[11][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][26] .is_wysiwyg = "true";
defparam \regs[11][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N17
dffeas \regs[10][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][26] .is_wysiwyg = "true";
defparam \regs[10][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N21
dffeas \regs[8][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][26] .is_wysiwyg = "true";
defparam \regs[8][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N20
cycloneive_lcell_comb \Mux37~10 (
// Equation(s):
// \Mux37~10_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][26]~q )) # (!dcifimemload_17 & ((\regs[8][26]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][26]~q ),
	.datac(\regs[8][26]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux37~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~10 .lut_mask = 16'hEE50;
defparam \Mux37~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N30
cycloneive_lcell_comb \Mux37~11 (
// Equation(s):
// \Mux37~11_combout  = (dcifimemload_16 & ((\Mux37~10_combout  & ((\regs[11][26]~q ))) # (!\Mux37~10_combout  & (\regs[9][26]~q )))) # (!dcifimemload_16 & (((\Mux37~10_combout ))))

	.dataa(\regs[9][26]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[11][26]~q ),
	.datad(\Mux37~10_combout ),
	.cin(gnd),
	.combout(\Mux37~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~11 .lut_mask = 16'hF388;
defparam \Mux37~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N27
dffeas \regs[14][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][26] .is_wysiwyg = "true";
defparam \regs[14][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N7
dffeas \regs[15][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][26] .is_wysiwyg = "true";
defparam \regs[15][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N29
dffeas \regs[12][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][26] .is_wysiwyg = "true";
defparam \regs[12][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N28
cycloneive_lcell_comb \Mux37~17 (
// Equation(s):
// \Mux37~17_combout  = (dcifimemload_16 & ((\regs[13][26]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[12][26]~q  & !dcifimemload_17))))

	.dataa(\regs[13][26]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[12][26]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux37~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~17 .lut_mask = 16'hCCB8;
defparam \Mux37~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N6
cycloneive_lcell_comb \Mux37~18 (
// Equation(s):
// \Mux37~18_combout  = (dcifimemload_17 & ((\Mux37~17_combout  & ((\regs[15][26]~q ))) # (!\Mux37~17_combout  & (\regs[14][26]~q )))) # (!dcifimemload_17 & (((\Mux37~17_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[14][26]~q ),
	.datac(\regs[15][26]~q ),
	.datad(\Mux37~17_combout ),
	.cin(gnd),
	.combout(\Mux37~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~18 .lut_mask = 16'hF588;
defparam \Mux37~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N9
dffeas \regs[6][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][26] .is_wysiwyg = "true";
defparam \regs[6][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N3
dffeas \regs[7][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][26] .is_wysiwyg = "true";
defparam \regs[7][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N25
dffeas \regs[4][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][26] .is_wysiwyg = "true";
defparam \regs[4][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N24
cycloneive_lcell_comb \Mux37~12 (
// Equation(s):
// \Mux37~12_combout  = (dcifimemload_16 & ((\regs[5][26]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][26]~q  & !dcifimemload_17))))

	.dataa(\regs[5][26]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][26]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux37~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~12 .lut_mask = 16'hCCB8;
defparam \Mux37~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N2
cycloneive_lcell_comb \Mux37~13 (
// Equation(s):
// \Mux37~13_combout  = (dcifimemload_17 & ((\Mux37~12_combout  & ((\regs[7][26]~q ))) # (!\Mux37~12_combout  & (\regs[6][26]~q )))) # (!dcifimemload_17 & (((\Mux37~12_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][26]~q ),
	.datac(\regs[7][26]~q ),
	.datad(\Mux37~12_combout ),
	.cin(gnd),
	.combout(\Mux37~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~13 .lut_mask = 16'hF588;
defparam \Mux37~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N7
dffeas \regs[2][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][26] .is_wysiwyg = "true";
defparam \regs[2][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N31
dffeas \regs[3][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][26] .is_wysiwyg = "true";
defparam \regs[3][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N1
dffeas \regs[1][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][26] .is_wysiwyg = "true";
defparam \regs[1][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N0
cycloneive_lcell_comb \Mux37~14 (
// Equation(s):
// \Mux37~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][26]~q )) # (!dcifimemload_17 & ((\regs[1][26]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[3][26]~q ),
	.datac(\regs[1][26]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux37~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~14 .lut_mask = 16'h88A0;
defparam \Mux37~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N6
cycloneive_lcell_comb \Mux37~15 (
// Equation(s):
// \Mux37~15_combout  = (\Mux37~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][26]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][26]~q ),
	.datad(\Mux37~14_combout ),
	.cin(gnd),
	.combout(\Mux37~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~15 .lut_mask = 16'hFF40;
defparam \Mux37~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N20
cycloneive_lcell_comb \Mux37~16 (
// Equation(s):
// \Mux37~16_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\Mux37~13_combout )) # (!dcifimemload_18 & ((\Mux37~15_combout )))))

	.dataa(\Mux37~13_combout ),
	.datab(dcifimemload_19),
	.datac(dcifimemload_18),
	.datad(\Mux37~15_combout ),
	.cin(gnd),
	.combout(\Mux37~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~16 .lut_mask = 16'hE3E0;
defparam \Mux37~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N10
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (dcifimemload_24 & (((\regs[27][26]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[19][26]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[19][26]~q ),
	.datac(\regs[27][26]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'hAAE4;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N16
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// \Mux5~8_combout  = (dcifimemload_23 & ((\Mux5~7_combout  & (\regs[31][26]~q )) # (!\Mux5~7_combout  & ((\regs[23][26]~q ))))) # (!dcifimemload_23 & (((\Mux5~7_combout ))))

	.dataa(\regs[31][26]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[23][26]~q ),
	.datad(\Mux5~7_combout ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hBBC0;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N8
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (dcifimemload_24 & (((\regs[25][26]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[17][26]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[17][26]~q ),
	.datac(\regs[25][26]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hAAE4;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N10
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (\Mux5~0_combout  & ((\regs[29][26]~q ) # ((!dcifimemload_23)))) # (!\Mux5~0_combout  & (((\regs[21][26]~q  & dcifimemload_23))))

	.dataa(\regs[29][26]~q ),
	.datab(\regs[21][26]~q ),
	.datac(\Mux5~0_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hACF0;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N27
dffeas \regs[26][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][26] .is_wysiwyg = "true";
defparam \regs[26][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N23
dffeas \regs[18][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][26] .is_wysiwyg = "true";
defparam \regs[18][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N6
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (dcifimemload_23 & (((\regs[22][26]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[18][26]~q  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[18][26]~q ),
	.datac(\regs[22][26]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hAAE4;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N26
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (dcifimemload_24 & ((\Mux5~2_combout  & (\regs[30][26]~q )) # (!\Mux5~2_combout  & ((\regs[26][26]~q ))))) # (!dcifimemload_24 & (((\Mux5~2_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[30][26]~q ),
	.datac(\regs[26][26]~q ),
	.datad(\Mux5~2_combout ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hDDA0;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N18
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[20][26]~q ))) # (!dcifimemload_23 & (\regs[16][26]~q ))))

	.dataa(dcifimemload_24),
	.datab(\regs[16][26]~q ),
	.datac(\regs[20][26]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hFA44;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N0
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (dcifimemload_24 & ((\Mux5~4_combout  & (\regs[28][26]~q )) # (!\Mux5~4_combout  & ((\regs[24][26]~q ))))) # (!dcifimemload_24 & (((\Mux5~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[28][26]~q ),
	.datac(\regs[24][26]~q ),
	.datad(\Mux5~4_combout ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hDDA0;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N0
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux5~3_combout )) # (!dcifimemload_22 & ((\Mux5~5_combout )))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux5~3_combout ),
	.datad(\Mux5~5_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hD9C8;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N26
cycloneive_lcell_comb \Mux5~9 (
// Equation(s):
// \Mux5~9_combout  = (dcifimemload_21 & ((\Mux5~6_combout  & (\Mux5~8_combout )) # (!\Mux5~6_combout  & ((\Mux5~1_combout ))))) # (!dcifimemload_21 & (((\Mux5~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux5~8_combout ),
	.datac(\Mux5~1_combout ),
	.datad(\Mux5~6_combout ),
	.cin(gnd),
	.combout(\Mux5~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~9 .lut_mask = 16'hDDA0;
defparam \Mux5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \Mux5~12 (
// Equation(s):
// \Mux5~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][26]~q ))) # (!dcifimemload_22 & (\regs[8][26]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][26]~q ),
	.datac(\regs[10][26]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux5~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~12 .lut_mask = 16'hFA44;
defparam \Mux5~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N8
cycloneive_lcell_comb \Mux5~13 (
// Equation(s):
// \Mux5~13_combout  = (dcifimemload_21 & ((\Mux5~12_combout  & (\regs[11][26]~q )) # (!\Mux5~12_combout  & ((\regs[9][26]~q ))))) # (!dcifimemload_21 & (((\Mux5~12_combout ))))

	.dataa(\regs[11][26]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[9][26]~q ),
	.datad(\Mux5~12_combout ),
	.cin(gnd),
	.combout(\Mux5~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~13 .lut_mask = 16'hBBC0;
defparam \Mux5~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N30
cycloneive_lcell_comb \Mux5~14 (
// Equation(s):
// \Mux5~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][26]~q ))) # (!dcifimemload_22 & (\regs[1][26]~q ))))

	.dataa(\regs[1][26]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[3][26]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux5~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~14 .lut_mask = 16'hC088;
defparam \Mux5~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N16
cycloneive_lcell_comb \Mux5~15 (
// Equation(s):
// \Mux5~15_combout  = (\Mux5~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \regs[2][26]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[2][26]~q ),
	.datad(\Mux5~14_combout ),
	.cin(gnd),
	.combout(\Mux5~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~15 .lut_mask = 16'hFF40;
defparam \Mux5~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N2
cycloneive_lcell_comb \Mux5~16 (
// Equation(s):
// \Mux5~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux5~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & ((\Mux5~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux5~13_combout ),
	.datad(\Mux5~15_combout ),
	.cin(gnd),
	.combout(\Mux5~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~16 .lut_mask = 16'hB9A8;
defparam \Mux5~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N17
dffeas \regs[13][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~16_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][26] .is_wysiwyg = "true";
defparam \regs[13][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N16
cycloneive_lcell_comb \Mux5~17 (
// Equation(s):
// \Mux5~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\regs[13][26]~q ))) # (!dcifimemload_21 & (\regs[12][26]~q ))))

	.dataa(\regs[12][26]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[13][26]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux5~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~17 .lut_mask = 16'hFC22;
defparam \Mux5~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N26
cycloneive_lcell_comb \Mux5~18 (
// Equation(s):
// \Mux5~18_combout  = (dcifimemload_22 & ((\Mux5~17_combout  & (\regs[15][26]~q )) # (!\Mux5~17_combout  & ((\regs[14][26]~q ))))) # (!dcifimemload_22 & (((\Mux5~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][26]~q ),
	.datac(\regs[14][26]~q ),
	.datad(\Mux5~17_combout ),
	.cin(gnd),
	.combout(\Mux5~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~18 .lut_mask = 16'hDDA0;
defparam \Mux5~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N8
cycloneive_lcell_comb \Mux5~11 (
// Equation(s):
// \Mux5~11_combout  = (\Mux5~10_combout  & (((\regs[7][26]~q )) # (!dcifimemload_22))) # (!\Mux5~10_combout  & (dcifimemload_22 & (\regs[6][26]~q )))

	.dataa(\Mux5~10_combout ),
	.datab(dcifimemload_22),
	.datac(\regs[6][26]~q ),
	.datad(\regs[7][26]~q ),
	.cin(gnd),
	.combout(\Mux5~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~11 .lut_mask = 16'hEA62;
defparam \Mux5~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N28
cycloneive_lcell_comb \Mux5~19 (
// Equation(s):
// \Mux5~19_combout  = (dcifimemload_23 & ((\Mux5~16_combout  & (\Mux5~18_combout )) # (!\Mux5~16_combout  & ((\Mux5~11_combout ))))) # (!dcifimemload_23 & (\Mux5~16_combout ))

	.dataa(dcifimemload_23),
	.datab(\Mux5~16_combout ),
	.datac(\Mux5~18_combout ),
	.datad(\Mux5~11_combout ),
	.cin(gnd),
	.combout(\Mux5~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~19 .lut_mask = 16'hE6C4;
defparam \Mux5~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N28
cycloneive_lcell_comb \regs~17 (
// Equation(s):
// \regs~17_combout  = (cuifRegSel_0 & ((cuifRegSel_11 & ((dcifimemload_9))) # (!cuifRegSel_11 & (ramiframload_25)))) # (!cuifRegSel_0 & (((cuifRegSel_11))))

	.dataa(ramiframload_25),
	.datab(cuifRegSel_0),
	.datac(dcifimemload_9),
	.datad(cuifRegSel_11),
	.cin(gnd),
	.combout(\regs~17_combout ),
	.cout());
// synopsys translate_off
defparam \regs~17 .lut_mask = 16'hF388;
defparam \regs~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N18
cycloneive_lcell_comb \regs~18 (
// Equation(s):
// \regs~18_combout  = (cuifRegSel_0) # ((\regs~17_combout  & (\Add1~46_combout )) # (!\regs~17_combout  & ((Selector0))))

	.dataa(Add115),
	.datab(cuifRegSel_0),
	.datac(\regs~17_combout ),
	.datad(Selector0),
	.cin(gnd),
	.combout(\regs~18_combout ),
	.cout());
// synopsys translate_off
defparam \regs~18 .lut_mask = 16'hEFEC;
defparam \regs~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N12
cycloneive_lcell_comb \regs~19 (
// Equation(s):
// \regs~19_combout  = (!\Equal0~1_combout  & ((\regs~17_combout  & (\regs~18_combout )) # (!\regs~17_combout  & (!\regs~18_combout  & Mux64))))

	.dataa(\regs~17_combout ),
	.datab(\regs~18_combout ),
	.datac(\Equal0~1_combout ),
	.datad(Mux64),
	.cin(gnd),
	.combout(\regs~19_combout ),
	.cout());
// synopsys translate_off
defparam \regs~19 .lut_mask = 16'h0908;
defparam \regs~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N27
dffeas \regs[28][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][25] .is_wysiwyg = "true";
defparam \regs[28][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N15
dffeas \regs[20][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][25] .is_wysiwyg = "true";
defparam \regs[20][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N17
dffeas \regs[16][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][25] .is_wysiwyg = "true";
defparam \regs[16][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N16
cycloneive_lcell_comb \Mux38~4 (
// Equation(s):
// \Mux38~4_combout  = (dcifimemload_18 & ((\regs[20][25]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[16][25]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[20][25]~q ),
	.datac(\regs[16][25]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux38~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~4 .lut_mask = 16'hAAD8;
defparam \Mux38~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N26
cycloneive_lcell_comb \Mux38~5 (
// Equation(s):
// \Mux38~5_combout  = (dcifimemload_19 & ((\Mux38~4_combout  & ((\regs[28][25]~q ))) # (!\Mux38~4_combout  & (\regs[24][25]~q )))) # (!dcifimemload_19 & (((\Mux38~4_combout ))))

	.dataa(\regs[24][25]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[28][25]~q ),
	.datad(\Mux38~4_combout ),
	.cin(gnd),
	.combout(\Mux38~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~5 .lut_mask = 16'hF388;
defparam \Mux38~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N29
dffeas \regs[30][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][25] .is_wysiwyg = "true";
defparam \regs[30][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N7
dffeas \regs[18][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][25] .is_wysiwyg = "true";
defparam \regs[18][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N6
cycloneive_lcell_comb \Mux38~2 (
// Equation(s):
// \Mux38~2_combout  = (dcifimemload_18 & ((\regs[22][25]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[18][25]~q  & !dcifimemload_19))))

	.dataa(\regs[22][25]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][25]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~2 .lut_mask = 16'hCCB8;
defparam \Mux38~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N28
cycloneive_lcell_comb \Mux38~3 (
// Equation(s):
// \Mux38~3_combout  = (dcifimemload_19 & ((\Mux38~2_combout  & ((\regs[30][25]~q ))) # (!\Mux38~2_combout  & (\regs[26][25]~q )))) # (!dcifimemload_19 & (((\Mux38~2_combout ))))

	.dataa(\regs[26][25]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[30][25]~q ),
	.datad(\Mux38~2_combout ),
	.cin(gnd),
	.combout(\Mux38~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~3 .lut_mask = 16'hF388;
defparam \Mux38~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N12
cycloneive_lcell_comb \Mux38~6 (
// Equation(s):
// \Mux38~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux38~3_combout ))) # (!dcifimemload_17 & (\Mux38~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux38~5_combout ),
	.datad(\Mux38~3_combout ),
	.cin(gnd),
	.combout(\Mux38~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~6 .lut_mask = 16'hDC98;
defparam \Mux38~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N8
cycloneive_lcell_comb \regs[21][25]~feeder (
// Equation(s):
// \regs[21][25]~feeder_combout  = \regs~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~19_combout ),
	.cin(gnd),
	.combout(\regs[21][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N9
dffeas \regs[21][25] (
	.clk(CLK),
	.d(\regs[21][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][25] .is_wysiwyg = "true";
defparam \regs[21][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N15
dffeas \regs[25][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][25] .is_wysiwyg = "true";
defparam \regs[25][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N29
dffeas \regs[17][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][25] .is_wysiwyg = "true";
defparam \regs[17][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N28
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[25][25]~q )) # (!dcifimemload_19 & ((\regs[17][25]~q )))))

	.dataa(dcifimemload_18),
	.datab(\regs[25][25]~q ),
	.datac(\regs[17][25]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hEE50;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N13
dffeas \regs[29][25] (
	.clk(CLK),
	.d(\regs~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][25] .is_wysiwyg = "true";
defparam \regs[29][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N14
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (dcifimemload_18 & ((\Mux38~0_combout  & ((\regs[29][25]~q ))) # (!\Mux38~0_combout  & (\regs[21][25]~q )))) # (!dcifimemload_18 & (((\Mux38~0_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[21][25]~q ),
	.datac(\Mux38~0_combout ),
	.datad(\regs[29][25]~q ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hF858;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N26
cycloneive_lcell_comb \regs[31][25]~feeder (
// Equation(s):
// \regs[31][25]~feeder_combout  = \regs~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~19_combout ),
	.cin(gnd),
	.combout(\regs[31][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[31][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N27
dffeas \regs[31][25] (
	.clk(CLK),
	.d(\regs[31][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][25] .is_wysiwyg = "true";
defparam \regs[31][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N19
dffeas \regs[23][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][25] .is_wysiwyg = "true";
defparam \regs[23][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N14
cycloneive_lcell_comb \regs[27][25]~feeder (
// Equation(s):
// \regs[27][25]~feeder_combout  = \regs~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~19_combout ),
	.cin(gnd),
	.combout(\regs[27][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N15
dffeas \regs[27][25] (
	.clk(CLK),
	.d(\regs[27][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][25] .is_wysiwyg = "true";
defparam \regs[27][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N20
cycloneive_lcell_comb \Mux38~7 (
// Equation(s):
// \Mux38~7_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[27][25]~q ))) # (!dcifimemload_19 & (\regs[19][25]~q ))))

	.dataa(\regs[19][25]~q ),
	.datab(\regs[27][25]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux38~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~7 .lut_mask = 16'hFC0A;
defparam \Mux38~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N28
cycloneive_lcell_comb \Mux38~8 (
// Equation(s):
// \Mux38~8_combout  = (dcifimemload_18 & ((\Mux38~7_combout  & (\regs[31][25]~q )) # (!\Mux38~7_combout  & ((\regs[23][25]~q ))))) # (!dcifimemload_18 & (((\Mux38~7_combout ))))

	.dataa(\regs[31][25]~q ),
	.datab(\regs[23][25]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux38~7_combout ),
	.cin(gnd),
	.combout(\Mux38~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~8 .lut_mask = 16'hAFC0;
defparam \Mux38~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N29
dffeas \regs[6][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][25] .is_wysiwyg = "true";
defparam \regs[6][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N29
dffeas \regs[4][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][25] .is_wysiwyg = "true";
defparam \regs[4][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N28
cycloneive_lcell_comb \Mux38~10 (
// Equation(s):
// \Mux38~10_combout  = (dcifimemload_16 & ((\regs[5][25]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][25]~q  & !dcifimemload_17))))

	.dataa(\regs[5][25]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][25]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux38~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~10 .lut_mask = 16'hCCB8;
defparam \Mux38~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N27
dffeas \regs[7][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][25] .is_wysiwyg = "true";
defparam \regs[7][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N26
cycloneive_lcell_comb \Mux38~11 (
// Equation(s):
// \Mux38~11_combout  = (\Mux38~10_combout  & (((\regs[7][25]~q ) # (!dcifimemload_17)))) # (!\Mux38~10_combout  & (\regs[6][25]~q  & ((dcifimemload_17))))

	.dataa(\regs[6][25]~q ),
	.datab(\Mux38~10_combout ),
	.datac(\regs[7][25]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux38~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~11 .lut_mask = 16'hE2CC;
defparam \Mux38~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N31
dffeas \regs[14][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][25] .is_wysiwyg = "true";
defparam \regs[14][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N15
dffeas \regs[15][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][25] .is_wysiwyg = "true";
defparam \regs[15][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N1
dffeas \regs[12][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][25] .is_wysiwyg = "true";
defparam \regs[12][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N0
cycloneive_lcell_comb \Mux38~17 (
// Equation(s):
// \Mux38~17_combout  = (dcifimemload_16 & ((\regs[13][25]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[12][25]~q  & !dcifimemload_17))))

	.dataa(\regs[13][25]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[12][25]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux38~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~17 .lut_mask = 16'hCCB8;
defparam \Mux38~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N14
cycloneive_lcell_comb \Mux38~18 (
// Equation(s):
// \Mux38~18_combout  = (dcifimemload_17 & ((\Mux38~17_combout  & ((\regs[15][25]~q ))) # (!\Mux38~17_combout  & (\regs[14][25]~q )))) # (!dcifimemload_17 & (((\Mux38~17_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[14][25]~q ),
	.datac(\regs[15][25]~q ),
	.datad(\Mux38~17_combout ),
	.cin(gnd),
	.combout(\Mux38~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~18 .lut_mask = 16'hF588;
defparam \Mux38~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N17
dffeas \regs[9][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][25] .is_wysiwyg = "true";
defparam \regs[9][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N19
dffeas \regs[11][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][25] .is_wysiwyg = "true";
defparam \regs[11][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N13
dffeas \regs[8][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][25] .is_wysiwyg = "true";
defparam \regs[8][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N12
cycloneive_lcell_comb \Mux38~12 (
// Equation(s):
// \Mux38~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][25]~q )) # (!dcifimemload_17 & ((\regs[8][25]~q )))))

	.dataa(\regs[10][25]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[8][25]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux38~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~12 .lut_mask = 16'hEE30;
defparam \Mux38~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N18
cycloneive_lcell_comb \Mux38~13 (
// Equation(s):
// \Mux38~13_combout  = (dcifimemload_16 & ((\Mux38~12_combout  & ((\regs[11][25]~q ))) # (!\Mux38~12_combout  & (\regs[9][25]~q )))) # (!dcifimemload_16 & (((\Mux38~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][25]~q ),
	.datac(\regs[11][25]~q ),
	.datad(\Mux38~12_combout ),
	.cin(gnd),
	.combout(\Mux38~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~13 .lut_mask = 16'hF588;
defparam \Mux38~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N24
cycloneive_lcell_comb \regs[3][25]~feeder (
// Equation(s):
// \regs[3][25]~feeder_combout  = \regs~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~19_combout ),
	.cin(gnd),
	.combout(\regs[3][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N25
dffeas \regs[3][25] (
	.clk(CLK),
	.d(\regs[3][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][25] .is_wysiwyg = "true";
defparam \regs[3][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N9
dffeas \regs[1][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][25] .is_wysiwyg = "true";
defparam \regs[1][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N8
cycloneive_lcell_comb \Mux38~14 (
// Equation(s):
// \Mux38~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][25]~q )) # (!dcifimemload_17 & ((\regs[1][25]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[3][25]~q ),
	.datac(\regs[1][25]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux38~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~14 .lut_mask = 16'h88A0;
defparam \Mux38~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N15
dffeas \regs[2][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][25] .is_wysiwyg = "true";
defparam \regs[2][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N14
cycloneive_lcell_comb \Mux38~15 (
// Equation(s):
// \Mux38~15_combout  = (\Mux38~14_combout ) # ((!dcifimemload_16 & (\regs[2][25]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\Mux38~14_combout ),
	.datac(\regs[2][25]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux38~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~15 .lut_mask = 16'hDCCC;
defparam \Mux38~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N20
cycloneive_lcell_comb \Mux38~16 (
// Equation(s):
// \Mux38~16_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & (\Mux38~13_combout )) # (!dcifimemload_19 & ((\Mux38~15_combout )))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux38~13_combout ),
	.datad(\Mux38~15_combout ),
	.cin(gnd),
	.combout(\Mux38~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~16 .lut_mask = 16'hD9C8;
defparam \Mux38~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N1
dffeas \regs[24][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][25] .is_wysiwyg = "true";
defparam \regs[24][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N0
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (dcifimemload_24 & (((\regs[24][25]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[16][25]~q  & ((!dcifimemload_23))))

	.dataa(\regs[16][25]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[24][25]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hCCE2;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N30
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (dcifimemload_23 & ((\Mux6~4_combout  & ((\regs[28][25]~q ))) # (!\Mux6~4_combout  & (\regs[20][25]~q )))) # (!dcifimemload_23 & (((\Mux6~4_combout ))))

	.dataa(\regs[20][25]~q ),
	.datab(\regs[28][25]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux6~4_combout ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'hCFA0;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N8
cycloneive_lcell_comb \regs[22][25]~feeder (
// Equation(s):
// \regs[22][25]~feeder_combout  = \regs~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~19_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[22][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][25]~feeder .lut_mask = 16'hF0F0;
defparam \regs[22][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N9
dffeas \regs[22][25] (
	.clk(CLK),
	.d(\regs[22][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][25] .is_wysiwyg = "true";
defparam \regs[22][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N1
dffeas \regs[26][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][25] .is_wysiwyg = "true";
defparam \regs[26][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N0
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\regs[26][25]~q ))) # (!dcifimemload_24 & (\regs[18][25]~q ))))

	.dataa(dcifimemload_23),
	.datab(\regs[18][25]~q ),
	.datac(\regs[26][25]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hFA44;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N28
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (\Mux6~2_combout  & ((\regs[30][25]~q ) # ((!dcifimemload_23)))) # (!\Mux6~2_combout  & (((\regs[22][25]~q  & dcifimemload_23))))

	.dataa(\regs[30][25]~q ),
	.datab(\regs[22][25]~q ),
	.datac(\Mux6~2_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hACF0;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N12
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux6~3_combout ))) # (!dcifimemload_22 & (\Mux6~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux6~5_combout ),
	.datad(\Mux6~3_combout ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hDC98;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N10
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[21][25]~q ))) # (!dcifimemload_23 & (\regs[17][25]~q ))))

	.dataa(\regs[17][25]~q ),
	.datab(\regs[21][25]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hFC0A;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N14
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (dcifimemload_24 & ((\Mux6~0_combout  & (\regs[29][25]~q )) # (!\Mux6~0_combout  & ((\regs[25][25]~q ))))) # (!dcifimemload_24 & (((\Mux6~0_combout ))))

	.dataa(\regs[29][25]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[25][25]~q ),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hBBC0;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N22
cycloneive_lcell_comb \regs[19][25]~feeder (
// Equation(s):
// \regs[19][25]~feeder_combout  = \regs~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~19_combout ),
	.cin(gnd),
	.combout(\regs[19][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[19][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N23
dffeas \regs[19][25] (
	.clk(CLK),
	.d(\regs[19][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][25] .is_wysiwyg = "true";
defparam \regs[19][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N18
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// \Mux6~7_combout  = (dcifimemload_23 & (((\regs[23][25]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[19][25]~q  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[19][25]~q ),
	.datac(\regs[23][25]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hAAE4;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N16
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (dcifimemload_24 & ((\Mux6~7_combout  & (\regs[31][25]~q )) # (!\Mux6~7_combout  & ((\regs[27][25]~q ))))) # (!dcifimemload_24 & (((\Mux6~7_combout ))))

	.dataa(\regs[31][25]~q ),
	.datab(\regs[27][25]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux6~7_combout ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'hAFC0;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N30
cycloneive_lcell_comb \Mux6~9 (
// Equation(s):
// \Mux6~9_combout  = (\Mux6~6_combout  & (((\Mux6~8_combout )) # (!dcifimemload_21))) # (!\Mux6~6_combout  & (dcifimemload_21 & (\Mux6~1_combout )))

	.dataa(\Mux6~6_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux6~1_combout ),
	.datad(\Mux6~8_combout ),
	.cin(gnd),
	.combout(\Mux6~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~9 .lut_mask = 16'hEA62;
defparam \Mux6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N30
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (\Mux6~17_combout  & ((\regs[15][25]~q ) # ((!dcifimemload_22)))) # (!\Mux6~17_combout  & (((\regs[14][25]~q  & dcifimemload_22))))

	.dataa(\Mux6~17_combout ),
	.datab(\regs[15][25]~q ),
	.datac(\regs[14][25]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hD8AA;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N5
dffeas \regs[10][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][25] .is_wysiwyg = "true";
defparam \regs[10][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N4
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][25]~q ))) # (!dcifimemload_22 & (\regs[8][25]~q ))))

	.dataa(\regs[8][25]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[10][25]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hFC22;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N22
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (\Mux6~10_combout  & ((\regs[11][25]~q ) # ((!dcifimemload_21)))) # (!\Mux6~10_combout  & (((\regs[9][25]~q  & dcifimemload_21))))

	.dataa(\regs[11][25]~q ),
	.datab(\regs[9][25]~q ),
	.datac(\Mux6~10_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hACF0;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N2
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][25]~q ))) # (!dcifimemload_22 & (\regs[1][25]~q ))))

	.dataa(\regs[1][25]~q ),
	.datab(\regs[3][25]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'hC0A0;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N4
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (\Mux6~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \regs[2][25]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[2][25]~q ),
	.datad(\Mux6~14_combout ),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'hFF40;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N11
dffeas \regs[5][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][25] .is_wysiwyg = "true";
defparam \regs[5][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N10
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (dcifimemload_21 & (((\regs[5][25]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][25]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][25]~q ),
	.datac(\regs[5][25]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hAAE4;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N28
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (dcifimemload_22 & ((\Mux6~12_combout  & (\regs[7][25]~q )) # (!\Mux6~12_combout  & ((\regs[6][25]~q ))))) # (!dcifimemload_22 & (((\Mux6~12_combout ))))

	.dataa(\regs[7][25]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[6][25]~q ),
	.datad(\Mux6~12_combout ),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hBBC0;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N18
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// \Mux6~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux6~13_combout ))) # (!dcifimemload_23 & (\Mux6~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux6~15_combout ),
	.datad(\Mux6~13_combout ),
	.cin(gnd),
	.combout(\Mux6~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hDC98;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N20
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// \Mux6~19_combout  = (dcifimemload_24 & ((\Mux6~16_combout  & (\Mux6~18_combout )) # (!\Mux6~16_combout  & ((\Mux6~11_combout ))))) # (!dcifimemload_24 & (((\Mux6~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux6~18_combout ),
	.datac(\Mux6~11_combout ),
	.datad(\Mux6~16_combout ),
	.cin(gnd),
	.combout(\Mux6~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'hDDA0;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N22
cycloneive_lcell_comb \regs~20 (
// Equation(s):
// \regs~20_combout  = (cuifRegSel_11 & ((cuifRegSel_0 & (dcifimemload_8)) # (!cuifRegSel_0 & ((\Add1~44_combout ))))) # (!cuifRegSel_11 & (((cuifRegSel_0))))

	.dataa(dcifimemload_8),
	.datab(Add114),
	.datac(cuifRegSel_11),
	.datad(cuifRegSel_0),
	.cin(gnd),
	.combout(\regs~20_combout ),
	.cout());
// synopsys translate_off
defparam \regs~20 .lut_mask = 16'hAFC0;
defparam \regs~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N28
cycloneive_lcell_comb \regs~21 (
// Equation(s):
// \regs~21_combout  = (cuifRegSel_11) # ((\regs~20_combout  & (ramiframload_24)) # (!\regs~20_combout  & ((Selector0))))

	.dataa(ramiframload_24),
	.datab(cuifRegSel_11),
	.datac(\regs~20_combout ),
	.datad(Selector0),
	.cin(gnd),
	.combout(\regs~21_combout ),
	.cout());
// synopsys translate_off
defparam \regs~21 .lut_mask = 16'hEFEC;
defparam \regs~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N6
cycloneive_lcell_comb \regs~22 (
// Equation(s):
// \regs~22_combout  = (!\Equal0~1_combout  & ((\regs~21_combout  & (\regs~20_combout )) # (!\regs~21_combout  & (!\regs~20_combout  & Mux71))))

	.dataa(\Equal0~1_combout ),
	.datab(\regs~21_combout ),
	.datac(\regs~20_combout ),
	.datad(Mux71),
	.cin(gnd),
	.combout(\regs~22_combout ),
	.cout());
// synopsys translate_off
defparam \regs~22 .lut_mask = 16'h4140;
defparam \regs~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N17
dffeas \regs[31][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][24] .is_wysiwyg = "true";
defparam \regs[31][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N23
dffeas \regs[27][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][24] .is_wysiwyg = "true";
defparam \regs[27][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N3
dffeas \regs[19][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][24] .is_wysiwyg = "true";
defparam \regs[19][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N25
dffeas \regs[23][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][24] .is_wysiwyg = "true";
defparam \regs[23][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N24
cycloneive_lcell_comb \Mux39~7 (
// Equation(s):
// \Mux39~7_combout  = (dcifimemload_18 & (((\regs[23][24]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[19][24]~q  & ((!dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[19][24]~q ),
	.datac(\regs[23][24]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux39~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~7 .lut_mask = 16'hAAE4;
defparam \Mux39~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N22
cycloneive_lcell_comb \Mux39~8 (
// Equation(s):
// \Mux39~8_combout  = (dcifimemload_19 & ((\Mux39~7_combout  & (\regs[31][24]~q )) # (!\Mux39~7_combout  & ((\regs[27][24]~q ))))) # (!dcifimemload_19 & (((\Mux39~7_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[31][24]~q ),
	.datac(\regs[27][24]~q ),
	.datad(\Mux39~7_combout ),
	.cin(gnd),
	.combout(\Mux39~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~8 .lut_mask = 16'hDDA0;
defparam \Mux39~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N13
dffeas \regs[29][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][24] .is_wysiwyg = "true";
defparam \regs[29][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N11
dffeas \regs[25][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][24] .is_wysiwyg = "true";
defparam \regs[25][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N3
dffeas \regs[21][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][24] .is_wysiwyg = "true";
defparam \regs[21][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N2
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (dcifimemload_18 & (((\regs[21][24]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[17][24]~q  & ((!dcifimemload_19))))

	.dataa(\regs[17][24]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[21][24]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hCCE2;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N10
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (dcifimemload_19 & ((\Mux39~0_combout  & (\regs[29][24]~q )) # (!\Mux39~0_combout  & ((\regs[25][24]~q ))))) # (!dcifimemload_19 & (((\Mux39~0_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[29][24]~q ),
	.datac(\regs[25][24]~q ),
	.datad(\Mux39~0_combout ),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hDDA0;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N27
dffeas \regs[28][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][24] .is_wysiwyg = "true";
defparam \regs[28][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N25
dffeas \regs[20][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][24] .is_wysiwyg = "true";
defparam \regs[20][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N24
cycloneive_lcell_comb \Mux39~5 (
// Equation(s):
// \Mux39~5_combout  = (\Mux39~4_combout  & ((\regs[28][24]~q ) # ((!dcifimemload_18)))) # (!\Mux39~4_combout  & (((\regs[20][24]~q  & dcifimemload_18))))

	.dataa(\Mux39~4_combout ),
	.datab(\regs[28][24]~q ),
	.datac(\regs[20][24]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux39~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~5 .lut_mask = 16'hD8AA;
defparam \Mux39~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y43_N13
dffeas \regs[22][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][24] .is_wysiwyg = "true";
defparam \regs[22][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y43_N11
dffeas \regs[26][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][24] .is_wysiwyg = "true";
defparam \regs[26][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N10
cycloneive_lcell_comb \Mux39~2 (
// Equation(s):
// \Mux39~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[26][24]~q ))) # (!dcifimemload_19 & (\regs[18][24]~q ))))

	.dataa(\regs[18][24]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[26][24]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux39~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~2 .lut_mask = 16'hFC22;
defparam \Mux39~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N12
cycloneive_lcell_comb \Mux39~3 (
// Equation(s):
// \Mux39~3_combout  = (dcifimemload_18 & ((\Mux39~2_combout  & (\regs[30][24]~q )) # (!\Mux39~2_combout  & ((\regs[22][24]~q ))))) # (!dcifimemload_18 & (((\Mux39~2_combout ))))

	.dataa(\regs[30][24]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[22][24]~q ),
	.datad(\Mux39~2_combout ),
	.cin(gnd),
	.combout(\Mux39~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~3 .lut_mask = 16'hBBC0;
defparam \Mux39~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N28
cycloneive_lcell_comb \Mux39~6 (
// Equation(s):
// \Mux39~6_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux39~3_combout ))) # (!dcifimemload_17 & (\Mux39~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux39~5_combout ),
	.datac(dcifimemload_17),
	.datad(\Mux39~3_combout ),
	.cin(gnd),
	.combout(\Mux39~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~6 .lut_mask = 16'hF4A4;
defparam \Mux39~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N12
cycloneive_lcell_comb \regs[14][24]~feeder (
// Equation(s):
// \regs[14][24]~feeder_combout  = \regs~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~22_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[14][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][24]~feeder .lut_mask = 16'hF0F0;
defparam \regs[14][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y44_N13
dffeas \regs[14][24] (
	.clk(CLK),
	.d(\regs[14][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][24] .is_wysiwyg = "true";
defparam \regs[14][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y44_N31
dffeas \regs[15][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][24] .is_wysiwyg = "true";
defparam \regs[15][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y44_N3
dffeas \regs[12][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][24] .is_wysiwyg = "true";
defparam \regs[12][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N2
cycloneive_lcell_comb \Mux39~17 (
// Equation(s):
// \Mux39~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][24]~q )) # (!dcifimemload_16 & ((\regs[12][24]~q )))))

	.dataa(\regs[13][24]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][24]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux39~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~17 .lut_mask = 16'hEE30;
defparam \Mux39~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N30
cycloneive_lcell_comb \Mux39~18 (
// Equation(s):
// \Mux39~18_combout  = (dcifimemload_17 & ((\Mux39~17_combout  & ((\regs[15][24]~q ))) # (!\Mux39~17_combout  & (\regs[14][24]~q )))) # (!dcifimemload_17 & (((\Mux39~17_combout ))))

	.dataa(\regs[14][24]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[15][24]~q ),
	.datad(\Mux39~17_combout ),
	.cin(gnd),
	.combout(\Mux39~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~18 .lut_mask = 16'hF388;
defparam \Mux39~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N27
dffeas \regs[10][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][24] .is_wysiwyg = "true";
defparam \regs[10][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N26
cycloneive_lcell_comb \Mux39~10 (
// Equation(s):
// \Mux39~10_combout  = (dcifimemload_17 & (((\regs[10][24]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\regs[8][24]~q  & ((!dcifimemload_16))))

	.dataa(\regs[8][24]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[10][24]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux39~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~10 .lut_mask = 16'hCCE2;
defparam \Mux39~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N31
dffeas \regs[11][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][24] .is_wysiwyg = "true";
defparam \regs[11][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N5
dffeas \regs[9][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][24] .is_wysiwyg = "true";
defparam \regs[9][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N4
cycloneive_lcell_comb \Mux39~11 (
// Equation(s):
// \Mux39~11_combout  = (\Mux39~10_combout  & ((\regs[11][24]~q ) # ((!dcifimemload_16)))) # (!\Mux39~10_combout  & (((\regs[9][24]~q  & dcifimemload_16))))

	.dataa(\Mux39~10_combout ),
	.datab(\regs[11][24]~q ),
	.datac(\regs[9][24]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux39~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~11 .lut_mask = 16'hD8AA;
defparam \Mux39~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N21
dffeas \regs[3][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][24] .is_wysiwyg = "true";
defparam \regs[3][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N1
dffeas \regs[1][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][24] .is_wysiwyg = "true";
defparam \regs[1][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N0
cycloneive_lcell_comb \Mux39~14 (
// Equation(s):
// \Mux39~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][24]~q )) # (!dcifimemload_17 & ((\regs[1][24]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[3][24]~q ),
	.datac(\regs[1][24]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux39~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~14 .lut_mask = 16'hD800;
defparam \Mux39~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N23
dffeas \regs[2][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][24] .is_wysiwyg = "true";
defparam \regs[2][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N22
cycloneive_lcell_comb \Mux39~15 (
// Equation(s):
// \Mux39~15_combout  = (\Mux39~14_combout ) # ((dcifimemload_17 & (\regs[2][24]~q  & !dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\Mux39~14_combout ),
	.datac(\regs[2][24]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux39~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~15 .lut_mask = 16'hCCEC;
defparam \Mux39~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N9
dffeas \regs[4][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][24] .is_wysiwyg = "true";
defparam \regs[4][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N8
cycloneive_lcell_comb \Mux39~12 (
// Equation(s):
// \Mux39~12_combout  = (dcifimemload_16 & ((\regs[5][24]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][24]~q  & !dcifimemload_17))))

	.dataa(\regs[5][24]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][24]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux39~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~12 .lut_mask = 16'hCCB8;
defparam \Mux39~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N7
dffeas \regs[7][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][24] .is_wysiwyg = "true";
defparam \regs[7][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N6
cycloneive_lcell_comb \Mux39~13 (
// Equation(s):
// \Mux39~13_combout  = (\Mux39~12_combout  & (((\regs[7][24]~q ) # (!dcifimemload_17)))) # (!\Mux39~12_combout  & (\regs[6][24]~q  & ((dcifimemload_17))))

	.dataa(\regs[6][24]~q ),
	.datab(\Mux39~12_combout ),
	.datac(\regs[7][24]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux39~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~13 .lut_mask = 16'hE2CC;
defparam \Mux39~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N16
cycloneive_lcell_comb \Mux39~16 (
// Equation(s):
// \Mux39~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux39~13_combout ))) # (!dcifimemload_18 & (\Mux39~15_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux39~15_combout ),
	.datad(\Mux39~13_combout ),
	.cin(gnd),
	.combout(\Mux39~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~16 .lut_mask = 16'hDC98;
defparam \Mux39~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N11
dffeas \regs[30][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][24] .is_wysiwyg = "true";
defparam \regs[30][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N10
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (\Mux7~2_combout  & (((\regs[30][24]~q ) # (!dcifimemload_24)))) # (!\Mux7~2_combout  & (\regs[26][24]~q  & ((dcifimemload_24))))

	.dataa(\Mux7~2_combout ),
	.datab(\regs[26][24]~q ),
	.datac(\regs[30][24]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hE4AA;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N29
dffeas \regs[16][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][24] .is_wysiwyg = "true";
defparam \regs[16][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N28
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (dcifimemload_23 & ((\regs[20][24]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[16][24]~q  & !dcifimemload_24))))

	.dataa(\regs[20][24]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[16][24]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'hCCB8;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N26
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (dcifimemload_24 & ((\Mux7~4_combout  & ((\regs[28][24]~q ))) # (!\Mux7~4_combout  & (\regs[24][24]~q )))) # (!dcifimemload_24 & (((\Mux7~4_combout ))))

	.dataa(\regs[24][24]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[28][24]~q ),
	.datad(\Mux7~4_combout ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hF388;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N4
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux7~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux7~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux7~3_combout ),
	.datad(\Mux7~5_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hB9A8;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N1
dffeas \regs[17][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][24] .is_wysiwyg = "true";
defparam \regs[17][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N0
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (dcifimemload_24 & ((\regs[25][24]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[17][24]~q  & !dcifimemload_23))))

	.dataa(\regs[25][24]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[17][24]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hCCB8;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N12
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (dcifimemload_23 & ((\Mux7~0_combout  & ((\regs[29][24]~q ))) # (!\Mux7~0_combout  & (\regs[21][24]~q )))) # (!dcifimemload_23 & (((\Mux7~0_combout ))))

	.dataa(\regs[21][24]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[29][24]~q ),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hF388;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N2
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (dcifimemload_24 & ((\regs[27][24]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[19][24]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][24]~q ),
	.datac(\regs[19][24]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hAAD8;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N16
cycloneive_lcell_comb \Mux7~8 (
// Equation(s):
// \Mux7~8_combout  = (dcifimemload_23 & ((\Mux7~7_combout  & ((\regs[31][24]~q ))) # (!\Mux7~7_combout  & (\regs[23][24]~q )))) # (!dcifimemload_23 & (((\Mux7~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[23][24]~q ),
	.datac(\regs[31][24]~q ),
	.datad(\Mux7~7_combout ),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~8 .lut_mask = 16'hF588;
defparam \Mux7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N14
cycloneive_lcell_comb \Mux7~9 (
// Equation(s):
// \Mux7~9_combout  = (dcifimemload_21 & ((\Mux7~6_combout  & ((\Mux7~8_combout ))) # (!\Mux7~6_combout  & (\Mux7~1_combout )))) # (!dcifimemload_21 & (\Mux7~6_combout ))

	.dataa(dcifimemload_21),
	.datab(\Mux7~6_combout ),
	.datac(\Mux7~1_combout ),
	.datad(\Mux7~8_combout ),
	.cin(gnd),
	.combout(\Mux7~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~9 .lut_mask = 16'hEC64;
defparam \Mux7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N8
cycloneive_lcell_comb \regs[6][24]~feeder (
// Equation(s):
// \regs[6][24]~feeder_combout  = \regs~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~22_combout ),
	.cin(gnd),
	.combout(\regs[6][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[6][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N9
dffeas \regs[6][24] (
	.clk(CLK),
	.d(\regs[6][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][24] .is_wysiwyg = "true";
defparam \regs[6][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N10
cycloneive_lcell_comb \Mux7~10 (
// Equation(s):
// \Mux7~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\regs[5][24]~q )) # (!dcifimemload_21 & ((\regs[4][24]~q )))))

	.dataa(\regs[5][24]~q ),
	.datab(\regs[4][24]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~10 .lut_mask = 16'hFA0C;
defparam \Mux7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N16
cycloneive_lcell_comb \Mux7~11 (
// Equation(s):
// \Mux7~11_combout  = (dcifimemload_22 & ((\Mux7~10_combout  & (\regs[7][24]~q )) # (!\Mux7~10_combout  & ((\regs[6][24]~q ))))) # (!dcifimemload_22 & (((\Mux7~10_combout ))))

	.dataa(\regs[7][24]~q ),
	.datab(\regs[6][24]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux7~10_combout ),
	.cin(gnd),
	.combout(\Mux7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~11 .lut_mask = 16'hAFC0;
defparam \Mux7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N12
cycloneive_lcell_comb \regs[13][24]~feeder (
// Equation(s):
// \regs[13][24]~feeder_combout  = \regs~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~22_combout ),
	.cin(gnd),
	.combout(\regs[13][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[13][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y44_N13
dffeas \regs[13][24] (
	.clk(CLK),
	.d(\regs[13][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][24] .is_wysiwyg = "true";
defparam \regs[13][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N30
cycloneive_lcell_comb \Mux7~17 (
// Equation(s):
// \Mux7~17_combout  = (dcifimemload_21 & ((\regs[13][24]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\regs[12][24]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[13][24]~q ),
	.datac(\regs[12][24]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux7~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~17 .lut_mask = 16'hAAD8;
defparam \Mux7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N24
cycloneive_lcell_comb \Mux7~18 (
// Equation(s):
// \Mux7~18_combout  = (\Mux7~17_combout  & (((\regs[15][24]~q ) # (!dcifimemload_22)))) # (!\Mux7~17_combout  & (\regs[14][24]~q  & ((dcifimemload_22))))

	.dataa(\regs[14][24]~q ),
	.datab(\regs[15][24]~q ),
	.datac(\Mux7~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~18 .lut_mask = 16'hCAF0;
defparam \Mux7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N25
dffeas \regs[8][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][24] .is_wysiwyg = "true";
defparam \regs[8][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N24
cycloneive_lcell_comb \Mux7~12 (
// Equation(s):
// \Mux7~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\regs[10][24]~q )) # (!dcifimemload_22 & ((\regs[8][24]~q )))))

	.dataa(\regs[10][24]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[8][24]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~12 .lut_mask = 16'hEE30;
defparam \Mux7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N30
cycloneive_lcell_comb \Mux7~13 (
// Equation(s):
// \Mux7~13_combout  = (dcifimemload_21 & ((\Mux7~12_combout  & ((\regs[11][24]~q ))) # (!\Mux7~12_combout  & (\regs[9][24]~q )))) # (!dcifimemload_21 & (((\Mux7~12_combout ))))

	.dataa(\regs[9][24]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[11][24]~q ),
	.datad(\Mux7~12_combout ),
	.cin(gnd),
	.combout(\Mux7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~13 .lut_mask = 16'hF388;
defparam \Mux7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N20
cycloneive_lcell_comb \Mux7~14 (
// Equation(s):
// \Mux7~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][24]~q ))) # (!dcifimemload_22 & (\regs[1][24]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[1][24]~q ),
	.datac(\regs[3][24]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~14 .lut_mask = 16'hA088;
defparam \Mux7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N16
cycloneive_lcell_comb \Mux7~15 (
// Equation(s):
// \Mux7~15_combout  = (\Mux7~14_combout ) # ((\regs[2][24]~q  & (!dcifimemload_21 & dcifimemload_22)))

	.dataa(\regs[2][24]~q ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\Mux7~14_combout ),
	.cin(gnd),
	.combout(\Mux7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~15 .lut_mask = 16'hFF20;
defparam \Mux7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N6
cycloneive_lcell_comb \Mux7~16 (
// Equation(s):
// \Mux7~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & (\Mux7~13_combout )) # (!dcifimemload_24 & ((\Mux7~15_combout )))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux7~13_combout ),
	.datad(\Mux7~15_combout ),
	.cin(gnd),
	.combout(\Mux7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~16 .lut_mask = 16'hD9C8;
defparam \Mux7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N28
cycloneive_lcell_comb \Mux7~19 (
// Equation(s):
// \Mux7~19_combout  = (dcifimemload_23 & ((\Mux7~16_combout  & ((\Mux7~18_combout ))) # (!\Mux7~16_combout  & (\Mux7~11_combout )))) # (!dcifimemload_23 & (((\Mux7~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux7~11_combout ),
	.datac(\Mux7~18_combout ),
	.datad(\Mux7~16_combout ),
	.cin(gnd),
	.combout(\Mux7~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~19 .lut_mask = 16'hF588;
defparam \Mux7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N4
cycloneive_lcell_comb \regs~23 (
// Equation(s):
// \regs~23_combout  = (\Selector8~1_combout  & !\Equal0~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector8),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\regs~23_combout ),
	.cout());
// synopsys translate_off
defparam \regs~23 .lut_mask = 16'h00F0;
defparam \regs~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N3
dffeas \regs[29][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][23] .is_wysiwyg = "true";
defparam \regs[29][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N14
cycloneive_lcell_comb \regs[21][23]~feeder (
// Equation(s):
// \regs[21][23]~feeder_combout  = \regs~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~23_combout ),
	.cin(gnd),
	.combout(\regs[21][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][23]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N15
dffeas \regs[21][23] (
	.clk(CLK),
	.d(\regs[21][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][23] .is_wysiwyg = "true";
defparam \regs[21][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N20
cycloneive_lcell_comb \regs[25][23]~feeder (
// Equation(s):
// \regs[25][23]~feeder_combout  = \regs~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~23_combout ),
	.cin(gnd),
	.combout(\regs[25][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[25][23]~feeder .lut_mask = 16'hFF00;
defparam \regs[25][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N21
dffeas \regs[25][23] (
	.clk(CLK),
	.d(\regs[25][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][23] .is_wysiwyg = "true";
defparam \regs[25][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N18
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[25][23]~q ))) # (!dcifimemload_19 & (\regs[17][23]~q ))))

	.dataa(\regs[17][23]~q ),
	.datab(\regs[25][23]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hFC0A;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N4
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (dcifimemload_18 & ((\Mux40~0_combout  & (\regs[29][23]~q )) # (!\Mux40~0_combout  & ((\regs[21][23]~q ))))) # (!dcifimemload_18 & (((\Mux40~0_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[29][23]~q ),
	.datac(\regs[21][23]~q ),
	.datad(\Mux40~0_combout ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hDDA0;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y43_N5
dffeas \regs[26][23] (
	.clk(CLK),
	.d(\regs~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][23] .is_wysiwyg = "true";
defparam \regs[26][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N25
dffeas \regs[18][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][23] .is_wysiwyg = "true";
defparam \regs[18][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N28
cycloneive_lcell_comb \Mux40~2 (
// Equation(s):
// \Mux40~2_combout  = (dcifimemload_18 & ((\regs[22][23]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[18][23]~q  & !dcifimemload_19))))

	.dataa(\regs[22][23]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][23]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~2 .lut_mask = 16'hCCB8;
defparam \Mux40~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N30
cycloneive_lcell_comb \Mux40~3 (
// Equation(s):
// \Mux40~3_combout  = (dcifimemload_19 & ((\Mux40~2_combout  & (\regs[30][23]~q )) # (!\Mux40~2_combout  & ((\regs[26][23]~q ))))) # (!dcifimemload_19 & (((\Mux40~2_combout ))))

	.dataa(\regs[30][23]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[26][23]~q ),
	.datad(\Mux40~2_combout ),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~3 .lut_mask = 16'hBBC0;
defparam \Mux40~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N1
dffeas \regs[24][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][23] .is_wysiwyg = "true";
defparam \regs[24][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N19
dffeas \regs[20][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][23] .is_wysiwyg = "true";
defparam \regs[20][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N18
cycloneive_lcell_comb \Mux40~4 (
// Equation(s):
// \Mux40~4_combout  = (dcifimemload_18 & (((\regs[20][23]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[16][23]~q  & ((!dcifimemload_19))))

	.dataa(\regs[16][23]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[20][23]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~4 .lut_mask = 16'hCCE2;
defparam \Mux40~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N0
cycloneive_lcell_comb \Mux40~5 (
// Equation(s):
// \Mux40~5_combout  = (dcifimemload_19 & ((\Mux40~4_combout  & (\regs[28][23]~q )) # (!\Mux40~4_combout  & ((\regs[24][23]~q ))))) # (!dcifimemload_19 & (((\Mux40~4_combout ))))

	.dataa(\regs[28][23]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[24][23]~q ),
	.datad(\Mux40~4_combout ),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~5 .lut_mask = 16'hBBC0;
defparam \Mux40~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N4
cycloneive_lcell_comb \Mux40~6 (
// Equation(s):
// \Mux40~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux40~3_combout )) # (!dcifimemload_17 & ((\Mux40~5_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux40~3_combout ),
	.datad(\Mux40~5_combout ),
	.cin(gnd),
	.combout(\Mux40~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~6 .lut_mask = 16'hD9C8;
defparam \Mux40~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N19
dffeas \regs[31][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][23] .is_wysiwyg = "true";
defparam \regs[31][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N4
cycloneive_lcell_comb \regs[23][23]~feeder (
// Equation(s):
// \regs[23][23]~feeder_combout  = \regs~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~23_combout ),
	.cin(gnd),
	.combout(\regs[23][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][23]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N5
dffeas \regs[23][23] (
	.clk(CLK),
	.d(\regs[23][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][23] .is_wysiwyg = "true";
defparam \regs[23][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N0
cycloneive_lcell_comb \regs[27][23]~feeder (
// Equation(s):
// \regs[27][23]~feeder_combout  = \regs~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~23_combout ),
	.cin(gnd),
	.combout(\regs[27][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][23]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N1
dffeas \regs[27][23] (
	.clk(CLK),
	.d(\regs[27][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][23] .is_wysiwyg = "true";
defparam \regs[27][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N6
cycloneive_lcell_comb \Mux40~7 (
// Equation(s):
// \Mux40~7_combout  = (dcifimemload_19 & (((\regs[27][23]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\regs[19][23]~q  & ((!dcifimemload_18))))

	.dataa(\regs[19][23]~q ),
	.datab(\regs[27][23]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux40~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~7 .lut_mask = 16'hF0CA;
defparam \Mux40~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N30
cycloneive_lcell_comb \Mux40~8 (
// Equation(s):
// \Mux40~8_combout  = (dcifimemload_18 & ((\Mux40~7_combout  & (\regs[31][23]~q )) # (!\Mux40~7_combout  & ((\regs[23][23]~q ))))) # (!dcifimemload_18 & (((\Mux40~7_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[31][23]~q ),
	.datac(\regs[23][23]~q ),
	.datad(\Mux40~7_combout ),
	.cin(gnd),
	.combout(\Mux40~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~8 .lut_mask = 16'hDDA0;
defparam \Mux40~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N31
dffeas \regs[7][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][23] .is_wysiwyg = "true";
defparam \regs[7][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N9
dffeas \regs[6][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][23] .is_wysiwyg = "true";
defparam \regs[6][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N7
dffeas \regs[5][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][23] .is_wysiwyg = "true";
defparam \regs[5][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N6
cycloneive_lcell_comb \Mux40~10 (
// Equation(s):
// \Mux40~10_combout  = (dcifimemload_16 & (((\regs[5][23]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][23]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][23]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[5][23]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux40~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~10 .lut_mask = 16'hCCE2;
defparam \Mux40~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N8
cycloneive_lcell_comb \Mux40~11 (
// Equation(s):
// \Mux40~11_combout  = (dcifimemload_17 & ((\Mux40~10_combout  & (\regs[7][23]~q )) # (!\Mux40~10_combout  & ((\regs[6][23]~q ))))) # (!dcifimemload_17 & (((\Mux40~10_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[7][23]~q ),
	.datac(\regs[6][23]~q ),
	.datad(\Mux40~10_combout ),
	.cin(gnd),
	.combout(\Mux40~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~11 .lut_mask = 16'hDDA0;
defparam \Mux40~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y45_N30
cycloneive_lcell_comb \regs[14][23]~feeder (
// Equation(s):
// \regs[14][23]~feeder_combout  = \regs~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~23_combout ),
	.cin(gnd),
	.combout(\regs[14][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][23]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y45_N31
dffeas \regs[14][23] (
	.clk(CLK),
	.d(\regs[14][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][23] .is_wysiwyg = "true";
defparam \regs[14][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y44_N29
dffeas \regs[15][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][23] .is_wysiwyg = "true";
defparam \regs[15][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y44_N23
dffeas \regs[12][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][23] .is_wysiwyg = "true";
defparam \regs[12][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N22
cycloneive_lcell_comb \Mux40~17 (
// Equation(s):
// \Mux40~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][23]~q )) # (!dcifimemload_16 & ((\regs[12][23]~q )))))

	.dataa(\regs[13][23]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][23]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux40~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~17 .lut_mask = 16'hEE30;
defparam \Mux40~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N28
cycloneive_lcell_comb \Mux40~18 (
// Equation(s):
// \Mux40~18_combout  = (dcifimemload_17 & ((\Mux40~17_combout  & ((\regs[15][23]~q ))) # (!\Mux40~17_combout  & (\regs[14][23]~q )))) # (!dcifimemload_17 & (((\Mux40~17_combout ))))

	.dataa(\regs[14][23]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[15][23]~q ),
	.datad(\Mux40~17_combout ),
	.cin(gnd),
	.combout(\Mux40~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~18 .lut_mask = 16'hF388;
defparam \Mux40~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y45_N11
dffeas \regs[2][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][23] .is_wysiwyg = "true";
defparam \regs[2][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y45_N29
dffeas \regs[1][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][23] .is_wysiwyg = "true";
defparam \regs[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N28
cycloneive_lcell_comb \Mux40~14 (
// Equation(s):
// \Mux40~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][23]~q )) # (!dcifimemload_17 & ((\regs[1][23]~q )))))

	.dataa(\regs[3][23]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[1][23]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux40~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~14 .lut_mask = 16'hB800;
defparam \Mux40~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N10
cycloneive_lcell_comb \Mux40~15 (
// Equation(s):
// \Mux40~15_combout  = (\Mux40~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][23]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][23]~q ),
	.datad(\Mux40~14_combout ),
	.cin(gnd),
	.combout(\Mux40~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~15 .lut_mask = 16'hFF40;
defparam \Mux40~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N5
dffeas \regs[8][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][23] .is_wysiwyg = "true";
defparam \regs[8][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N4
cycloneive_lcell_comb \Mux40~12 (
// Equation(s):
// \Mux40~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][23]~q )) # (!dcifimemload_17 & ((\regs[8][23]~q )))))

	.dataa(\regs[10][23]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[8][23]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux40~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~12 .lut_mask = 16'hEE30;
defparam \Mux40~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N23
dffeas \regs[11][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][23] .is_wysiwyg = "true";
defparam \regs[11][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N19
dffeas \regs[9][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][23] .is_wysiwyg = "true";
defparam \regs[9][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N22
cycloneive_lcell_comb \Mux40~13 (
// Equation(s):
// \Mux40~13_combout  = (dcifimemload_16 & ((\Mux40~12_combout  & (\regs[11][23]~q )) # (!\Mux40~12_combout  & ((\regs[9][23]~q ))))) # (!dcifimemload_16 & (\Mux40~12_combout ))

	.dataa(dcifimemload_16),
	.datab(\Mux40~12_combout ),
	.datac(\regs[11][23]~q ),
	.datad(\regs[9][23]~q ),
	.cin(gnd),
	.combout(\Mux40~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~13 .lut_mask = 16'hE6C4;
defparam \Mux40~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N20
cycloneive_lcell_comb \Mux40~16 (
// Equation(s):
// \Mux40~16_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & ((\Mux40~13_combout ))) # (!dcifimemload_19 & (\Mux40~15_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux40~15_combout ),
	.datad(\Mux40~13_combout ),
	.cin(gnd),
	.combout(\Mux40~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~16 .lut_mask = 16'hDC98;
defparam \Mux40~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N22
cycloneive_lcell_comb \regs[22][23]~feeder (
// Equation(s):
// \regs[22][23]~feeder_combout  = \regs~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~23_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[22][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][23]~feeder .lut_mask = 16'hF0F0;
defparam \regs[22][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y43_N23
dffeas \regs[22][23] (
	.clk(CLK),
	.d(\regs[22][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][23] .is_wysiwyg = "true";
defparam \regs[22][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N3
dffeas \regs[30][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][23] .is_wysiwyg = "true";
defparam \regs[30][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N24
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[26][23]~q )) # (!dcifimemload_24 & ((\regs[18][23]~q )))))

	.dataa(\regs[26][23]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[18][23]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hEE30;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N2
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (dcifimemload_23 & ((\Mux8~2_combout  & ((\regs[30][23]~q ))) # (!\Mux8~2_combout  & (\regs[22][23]~q )))) # (!dcifimemload_23 & (((\Mux8~2_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[22][23]~q ),
	.datac(\regs[30][23]~q ),
	.datad(\Mux8~2_combout ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hF588;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N12
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (dcifimemload_22 & (((dcifimemload_21) # (\Mux8~3_combout )))) # (!dcifimemload_22 & (\Mux8~5_combout  & (!dcifimemload_21)))

	.dataa(\Mux8~5_combout ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux8~3_combout ),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hCEC2;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N17
dffeas \regs[19][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][23] .is_wysiwyg = "true";
defparam \regs[19][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N16
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[23][23]~q )) # (!dcifimemload_23 & ((\regs[19][23]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[23][23]~q ),
	.datac(\regs[19][23]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hEE50;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N18
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// \Mux8~8_combout  = (dcifimemload_24 & ((\Mux8~7_combout  & ((\regs[31][23]~q ))) # (!\Mux8~7_combout  & (\regs[27][23]~q )))) # (!dcifimemload_24 & (((\Mux8~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][23]~q ),
	.datac(\regs[31][23]~q ),
	.datad(\Mux8~7_combout ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hF588;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N17
dffeas \regs[17][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][23] .is_wysiwyg = "true";
defparam \regs[17][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N16
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[21][23]~q )) # (!dcifimemload_23 & ((\regs[17][23]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[21][23]~q ),
	.datac(\regs[17][23]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hEE50;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N2
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (dcifimemload_24 & ((\Mux8~0_combout  & ((\regs[29][23]~q ))) # (!\Mux8~0_combout  & (\regs[25][23]~q )))) # (!dcifimemload_24 & (((\Mux8~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[25][23]~q ),
	.datac(\regs[29][23]~q ),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hF588;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N26
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// \Mux8~9_combout  = (\Mux8~6_combout  & (((\Mux8~8_combout )) # (!dcifimemload_21))) # (!\Mux8~6_combout  & (dcifimemload_21 & ((\Mux8~1_combout ))))

	.dataa(\Mux8~6_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux8~8_combout ),
	.datad(\Mux8~1_combout ),
	.cin(gnd),
	.combout(\Mux8~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'hE6A2;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N8
cycloneive_lcell_comb \regs[13][23]~feeder (
// Equation(s):
// \regs[13][23]~feeder_combout  = \regs~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~23_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[13][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][23]~feeder .lut_mask = 16'hF0F0;
defparam \regs[13][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y44_N9
dffeas \regs[13][23] (
	.clk(CLK),
	.d(\regs[13][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][23] .is_wysiwyg = "true";
defparam \regs[13][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y45_N26
cycloneive_lcell_comb \Mux8~17 (
// Equation(s):
// \Mux8~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\regs[13][23]~q )) # (!dcifimemload_21 & ((\regs[12][23]~q )))))

	.dataa(dcifimemload_22),
	.datab(\regs[13][23]~q ),
	.datac(\regs[12][23]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux8~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~17 .lut_mask = 16'hEE50;
defparam \Mux8~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y45_N24
cycloneive_lcell_comb \Mux8~18 (
// Equation(s):
// \Mux8~18_combout  = (\Mux8~17_combout  & (((\regs[15][23]~q ) # (!dcifimemload_22)))) # (!\Mux8~17_combout  & (\regs[14][23]~q  & ((dcifimemload_22))))

	.dataa(\regs[14][23]~q ),
	.datab(\regs[15][23]~q ),
	.datac(\Mux8~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux8~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~18 .lut_mask = 16'hCAF0;
defparam \Mux8~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N29
dffeas \regs[10][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][23] .is_wysiwyg = "true";
defparam \regs[10][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N28
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\regs[10][23]~q )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\regs[8][23]~q ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[10][23]~q ),
	.datad(\regs[8][23]~q ),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hB9A8;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N18
cycloneive_lcell_comb \Mux8~11 (
// Equation(s):
// \Mux8~11_combout  = (dcifimemload_21 & ((\Mux8~10_combout  & (\regs[11][23]~q )) # (!\Mux8~10_combout  & ((\regs[9][23]~q ))))) # (!dcifimemload_21 & (((\Mux8~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\regs[11][23]~q ),
	.datac(\regs[9][23]~q ),
	.datad(\Mux8~10_combout ),
	.cin(gnd),
	.combout(\Mux8~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~11 .lut_mask = 16'hDDA0;
defparam \Mux8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y45_N8
cycloneive_lcell_comb \regs[3][23]~feeder (
// Equation(s):
// \regs[3][23]~feeder_combout  = \regs~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~23_combout ),
	.cin(gnd),
	.combout(\regs[3][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][23]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y45_N9
dffeas \regs[3][23] (
	.clk(CLK),
	.d(\regs[3][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][23] .is_wysiwyg = "true";
defparam \regs[3][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y45_N16
cycloneive_lcell_comb \Mux8~14 (
// Equation(s):
// \Mux8~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][23]~q ))) # (!dcifimemload_22 & (\regs[1][23]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[1][23]~q ),
	.datac(\regs[3][23]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux8~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~14 .lut_mask = 16'hA088;
defparam \Mux8~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N8
cycloneive_lcell_comb \Mux8~15 (
// Equation(s):
// \Mux8~15_combout  = (\Mux8~14_combout ) # ((\regs[2][23]~q  & (!dcifimemload_21 & dcifimemload_22)))

	.dataa(\regs[2][23]~q ),
	.datab(dcifimemload_21),
	.datac(\Mux8~14_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux8~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~15 .lut_mask = 16'hF2F0;
defparam \Mux8~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N25
dffeas \regs[4][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][23] .is_wysiwyg = "true";
defparam \regs[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N24
cycloneive_lcell_comb \Mux8~12 (
// Equation(s):
// \Mux8~12_combout  = (dcifimemload_21 & ((dcifimemload_22) # ((\regs[5][23]~q )))) # (!dcifimemload_21 & (!dcifimemload_22 & (\regs[4][23]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[4][23]~q ),
	.datad(\regs[5][23]~q ),
	.cin(gnd),
	.combout(\Mux8~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~12 .lut_mask = 16'hBA98;
defparam \Mux8~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N30
cycloneive_lcell_comb \Mux8~13 (
// Equation(s):
// \Mux8~13_combout  = (dcifimemload_22 & ((\Mux8~12_combout  & ((\regs[7][23]~q ))) # (!\Mux8~12_combout  & (\regs[6][23]~q )))) # (!dcifimemload_22 & (((\Mux8~12_combout ))))

	.dataa(\regs[6][23]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[7][23]~q ),
	.datad(\Mux8~12_combout ),
	.cin(gnd),
	.combout(\Mux8~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~13 .lut_mask = 16'hF388;
defparam \Mux8~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N2
cycloneive_lcell_comb \Mux8~16 (
// Equation(s):
// \Mux8~16_combout  = (dcifimemload_23 & (((\Mux8~13_combout ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\Mux8~15_combout  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\Mux8~15_combout ),
	.datac(\Mux8~13_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux8~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~16 .lut_mask = 16'hAAE4;
defparam \Mux8~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N0
cycloneive_lcell_comb \Mux8~19 (
// Equation(s):
// \Mux8~19_combout  = (dcifimemload_24 & ((\Mux8~16_combout  & (\Mux8~18_combout )) # (!\Mux8~16_combout  & ((\Mux8~11_combout ))))) # (!dcifimemload_24 & (((\Mux8~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux8~18_combout ),
	.datac(\Mux8~11_combout ),
	.datad(\Mux8~16_combout ),
	.cin(gnd),
	.combout(\Mux8~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~19 .lut_mask = 16'hDDA0;
defparam \Mux8~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N18
cycloneive_lcell_comb \regs~24 (
// Equation(s):
// \regs~24_combout  = (!\Equal0~1_combout  & \Selector9~1_combout )

	.dataa(gnd),
	.datab(\Equal0~1_combout ),
	.datac(gnd),
	.datad(Selector9),
	.cin(gnd),
	.combout(\regs~24_combout ),
	.cout());
// synopsys translate_off
defparam \regs~24 .lut_mask = 16'h3300;
defparam \regs~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N4
cycloneive_lcell_comb \regs[29][22]~feeder (
// Equation(s):
// \regs[29][22]~feeder_combout  = \regs~24_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~24_combout ),
	.cin(gnd),
	.combout(\regs[29][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][22]~feeder .lut_mask = 16'hFF00;
defparam \regs[29][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N5
dffeas \regs[29][22] (
	.clk(CLK),
	.d(\regs[29][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][22] .is_wysiwyg = "true";
defparam \regs[29][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N7
dffeas \regs[25][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][22] .is_wysiwyg = "true";
defparam \regs[25][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N15
dffeas \regs[21][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][22] .is_wysiwyg = "true";
defparam \regs[21][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N14
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (dcifimemload_18 & (((\regs[21][22]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[17][22]~q  & ((!dcifimemload_19))))

	.dataa(\regs[17][22]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[21][22]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hCCE2;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N6
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (dcifimemload_19 & ((\Mux41~0_combout  & (\regs[29][22]~q )) # (!\Mux41~0_combout  & ((\regs[25][22]~q ))))) # (!dcifimemload_19 & (((\Mux41~0_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[29][22]~q ),
	.datac(\regs[25][22]~q ),
	.datad(\Mux41~0_combout ),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hDDA0;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N4
cycloneive_lcell_comb \regs[27][22]~feeder (
// Equation(s):
// \regs[27][22]~feeder_combout  = \regs~24_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~24_combout ),
	.cin(gnd),
	.combout(\regs[27][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][22]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N5
dffeas \regs[27][22] (
	.clk(CLK),
	.d(\regs[27][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][22] .is_wysiwyg = "true";
defparam \regs[27][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N31
dffeas \regs[31][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][22] .is_wysiwyg = "true";
defparam \regs[31][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N4
cycloneive_lcell_comb \regs[23][22]~feeder (
// Equation(s):
// \regs[23][22]~feeder_combout  = \regs~24_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~24_combout ),
	.cin(gnd),
	.combout(\regs[23][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][22]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N5
dffeas \regs[23][22] (
	.clk(CLK),
	.d(\regs[23][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][22] .is_wysiwyg = "true";
defparam \regs[23][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N6
cycloneive_lcell_comb \Mux41~7 (
// Equation(s):
// \Mux41~7_combout  = (dcifimemload_18 & (((\regs[23][22]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[19][22]~q  & ((!dcifimemload_19))))

	.dataa(\regs[19][22]~q ),
	.datab(\regs[23][22]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux41~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~7 .lut_mask = 16'hF0CA;
defparam \Mux41~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N22
cycloneive_lcell_comb \Mux41~8 (
// Equation(s):
// \Mux41~8_combout  = (dcifimemload_19 & ((\Mux41~7_combout  & ((\regs[31][22]~q ))) # (!\Mux41~7_combout  & (\regs[27][22]~q )))) # (!dcifimemload_19 & (((\Mux41~7_combout ))))

	.dataa(\regs[27][22]~q ),
	.datab(\regs[31][22]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux41~7_combout ),
	.cin(gnd),
	.combout(\Mux41~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~8 .lut_mask = 16'hCFA0;
defparam \Mux41~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N31
dffeas \regs[28][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][22] .is_wysiwyg = "true";
defparam \regs[28][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N17
dffeas \regs[20][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][22] .is_wysiwyg = "true";
defparam \regs[20][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N11
dffeas \regs[24][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][22] .is_wysiwyg = "true";
defparam \regs[24][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N10
cycloneive_lcell_comb \Mux41~4 (
// Equation(s):
// \Mux41~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[24][22]~q ))) # (!dcifimemload_19 & (\regs[16][22]~q ))))

	.dataa(\regs[16][22]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[24][22]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~4 .lut_mask = 16'hFC22;
defparam \Mux41~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N16
cycloneive_lcell_comb \Mux41~5 (
// Equation(s):
// \Mux41~5_combout  = (dcifimemload_18 & ((\Mux41~4_combout  & (\regs[28][22]~q )) # (!\Mux41~4_combout  & ((\regs[20][22]~q ))))) # (!dcifimemload_18 & (((\Mux41~4_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[28][22]~q ),
	.datac(\regs[20][22]~q ),
	.datad(\Mux41~4_combout ),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~5 .lut_mask = 16'hDDA0;
defparam \Mux41~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N8
cycloneive_lcell_comb \regs[22][22]~feeder (
// Equation(s):
// \regs[22][22]~feeder_combout  = \regs~24_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~24_combout ),
	.cin(gnd),
	.combout(\regs[22][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][22]~feeder .lut_mask = 16'hFF00;
defparam \regs[22][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y43_N9
dffeas \regs[22][22] (
	.clk(CLK),
	.d(\regs[22][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][22] .is_wysiwyg = "true";
defparam \regs[22][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y43_N19
dffeas \regs[26][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][22] .is_wysiwyg = "true";
defparam \regs[26][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N18
cycloneive_lcell_comb \Mux41~2 (
// Equation(s):
// \Mux41~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[26][22]~q ))) # (!dcifimemload_19 & (\regs[18][22]~q ))))

	.dataa(\regs[18][22]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[26][22]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~2 .lut_mask = 16'hFC22;
defparam \Mux41~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N20
cycloneive_lcell_comb \Mux41~3 (
// Equation(s):
// \Mux41~3_combout  = (dcifimemload_18 & ((\Mux41~2_combout  & (\regs[30][22]~q )) # (!\Mux41~2_combout  & ((\regs[22][22]~q ))))) # (!dcifimemload_18 & (((\Mux41~2_combout ))))

	.dataa(\regs[30][22]~q ),
	.datab(\regs[22][22]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux41~2_combout ),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~3 .lut_mask = 16'hAFC0;
defparam \Mux41~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N16
cycloneive_lcell_comb \Mux41~6 (
// Equation(s):
// \Mux41~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux41~3_combout ))) # (!dcifimemload_17 & (\Mux41~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux41~5_combout ),
	.datad(\Mux41~3_combout ),
	.cin(gnd),
	.combout(\Mux41~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~6 .lut_mask = 16'hDC98;
defparam \Mux41~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N27
dffeas \regs[11][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][22] .is_wysiwyg = "true";
defparam \regs[11][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N17
dffeas \regs[9][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][22] .is_wysiwyg = "true";
defparam \regs[9][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N3
dffeas \regs[10][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][22] .is_wysiwyg = "true";
defparam \regs[10][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N2
cycloneive_lcell_comb \Mux41~10 (
// Equation(s):
// \Mux41~10_combout  = (dcifimemload_17 & (((\regs[10][22]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\regs[8][22]~q  & ((!dcifimemload_16))))

	.dataa(\regs[8][22]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[10][22]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux41~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~10 .lut_mask = 16'hCCE2;
defparam \Mux41~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N16
cycloneive_lcell_comb \Mux41~11 (
// Equation(s):
// \Mux41~11_combout  = (dcifimemload_16 & ((\Mux41~10_combout  & (\regs[11][22]~q )) # (!\Mux41~10_combout  & ((\regs[9][22]~q ))))) # (!dcifimemload_16 & (((\Mux41~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[11][22]~q ),
	.datac(\regs[9][22]~q ),
	.datad(\Mux41~10_combout ),
	.cin(gnd),
	.combout(\Mux41~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~11 .lut_mask = 16'hDDA0;
defparam \Mux41~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N31
dffeas \regs[7][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][22] .is_wysiwyg = "true";
defparam \regs[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N1
dffeas \regs[4][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][22] .is_wysiwyg = "true";
defparam \regs[4][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N0
cycloneive_lcell_comb \Mux41~12 (
// Equation(s):
// \Mux41~12_combout  = (dcifimemload_16 & ((\regs[5][22]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][22]~q  & !dcifimemload_17))))

	.dataa(\regs[5][22]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][22]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux41~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~12 .lut_mask = 16'hCCB8;
defparam \Mux41~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N30
cycloneive_lcell_comb \Mux41~13 (
// Equation(s):
// \Mux41~13_combout  = (dcifimemload_17 & ((\Mux41~12_combout  & ((\regs[7][22]~q ))) # (!\Mux41~12_combout  & (\regs[6][22]~q )))) # (!dcifimemload_17 & (((\Mux41~12_combout ))))

	.dataa(\regs[6][22]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[7][22]~q ),
	.datad(\Mux41~12_combout ),
	.cin(gnd),
	.combout(\Mux41~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~13 .lut_mask = 16'hF388;
defparam \Mux41~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y45_N23
dffeas \regs[2][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][22] .is_wysiwyg = "true";
defparam \regs[2][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y45_N21
dffeas \regs[1][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][22] .is_wysiwyg = "true";
defparam \regs[1][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N20
cycloneive_lcell_comb \Mux41~14 (
// Equation(s):
// \Mux41~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][22]~q )) # (!dcifimemload_17 & ((\regs[1][22]~q )))))

	.dataa(\regs[3][22]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][22]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux41~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~14 .lut_mask = 16'h88C0;
defparam \Mux41~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N22
cycloneive_lcell_comb \Mux41~15 (
// Equation(s):
// \Mux41~15_combout  = (\Mux41~14_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][22]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[2][22]~q ),
	.datad(\Mux41~14_combout ),
	.cin(gnd),
	.combout(\Mux41~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~15 .lut_mask = 16'hFF20;
defparam \Mux41~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N4
cycloneive_lcell_comb \Mux41~16 (
// Equation(s):
// \Mux41~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & (\Mux41~13_combout )) # (!dcifimemload_18 & ((\Mux41~15_combout )))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux41~13_combout ),
	.datad(\Mux41~15_combout ),
	.cin(gnd),
	.combout(\Mux41~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~16 .lut_mask = 16'hD9C8;
defparam \Mux41~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N26
cycloneive_lcell_comb \regs[14][22]~feeder (
// Equation(s):
// \regs[14][22]~feeder_combout  = \regs~24_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~24_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[14][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][22]~feeder .lut_mask = 16'hF0F0;
defparam \regs[14][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y44_N27
dffeas \regs[14][22] (
	.clk(CLK),
	.d(\regs[14][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][22] .is_wysiwyg = "true";
defparam \regs[14][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N8
cycloneive_lcell_comb \regs[15][22]~feeder (
// Equation(s):
// \regs[15][22]~feeder_combout  = \regs~24_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~24_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[15][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][22]~feeder .lut_mask = 16'hF0F0;
defparam \regs[15][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y44_N9
dffeas \regs[15][22] (
	.clk(CLK),
	.d(\regs[15][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][22] .is_wysiwyg = "true";
defparam \regs[15][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y43_N1
dffeas \regs[12][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][22] .is_wysiwyg = "true";
defparam \regs[12][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N0
cycloneive_lcell_comb \Mux41~17 (
// Equation(s):
// \Mux41~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][22]~q )) # (!dcifimemload_16 & ((\regs[12][22]~q )))))

	.dataa(\regs[13][22]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][22]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux41~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~17 .lut_mask = 16'hEE30;
defparam \Mux41~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N22
cycloneive_lcell_comb \Mux41~18 (
// Equation(s):
// \Mux41~18_combout  = (dcifimemload_17 & ((\Mux41~17_combout  & ((\regs[15][22]~q ))) # (!\Mux41~17_combout  & (\regs[14][22]~q )))) # (!dcifimemload_17 & (((\Mux41~17_combout ))))

	.dataa(\regs[14][22]~q ),
	.datab(\regs[15][22]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux41~17_combout ),
	.cin(gnd),
	.combout(\Mux41~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~18 .lut_mask = 16'hCFA0;
defparam \Mux41~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N23
dffeas \regs[30][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][22] .is_wysiwyg = "true";
defparam \regs[30][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N1
dffeas \regs[18][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][22] .is_wysiwyg = "true";
defparam \regs[18][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N0
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (dcifimemload_23 & ((\regs[22][22]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[18][22]~q  & !dcifimemload_24))))

	.dataa(\regs[22][22]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[18][22]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hCCB8;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N22
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (dcifimemload_24 & ((\Mux9~2_combout  & ((\regs[30][22]~q ))) # (!\Mux9~2_combout  & (\regs[26][22]~q )))) # (!dcifimemload_24 & (((\Mux9~2_combout ))))

	.dataa(\regs[26][22]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[30][22]~q ),
	.datad(\Mux9~2_combout ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hF388;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N12
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux9~3_combout ))) # (!dcifimemload_22 & (\Mux9~5_combout ))))

	.dataa(\Mux9~5_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux9~3_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hFC22;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N25
dffeas \regs[17][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][22] .is_wysiwyg = "true";
defparam \regs[17][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N24
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (dcifimemload_24 & ((\regs[25][22]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[17][22]~q  & !dcifimemload_23))))

	.dataa(\regs[25][22]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[17][22]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hCCB8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N6
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (dcifimemload_23 & ((\Mux9~0_combout  & ((\regs[29][22]~q ))) # (!\Mux9~0_combout  & (\regs[21][22]~q )))) # (!dcifimemload_23 & (((\Mux9~0_combout ))))

	.dataa(\regs[21][22]~q ),
	.datab(\regs[29][22]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hCFA0;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N21
dffeas \regs[19][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][22] .is_wysiwyg = "true";
defparam \regs[19][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N20
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// \Mux9~7_combout  = (dcifimemload_24 & ((\regs[27][22]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[19][22]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][22]~q ),
	.datac(\regs[19][22]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'hAAD8;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N30
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (dcifimemload_23 & ((\Mux9~7_combout  & ((\regs[31][22]~q ))) # (!\Mux9~7_combout  & (\regs[23][22]~q )))) # (!dcifimemload_23 & (((\Mux9~7_combout ))))

	.dataa(\regs[23][22]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[31][22]~q ),
	.datad(\Mux9~7_combout ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hF388;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N4
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// \Mux9~9_combout  = (dcifimemload_21 & ((\Mux9~6_combout  & ((\Mux9~8_combout ))) # (!\Mux9~6_combout  & (\Mux9~1_combout )))) # (!dcifimemload_21 & (\Mux9~6_combout ))

	.dataa(dcifimemload_21),
	.datab(\Mux9~6_combout ),
	.datac(\Mux9~1_combout ),
	.datad(\Mux9~8_combout ),
	.cin(gnd),
	.combout(\Mux9~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hEC64;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N1
dffeas \regs[6][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][22] .is_wysiwyg = "true";
defparam \regs[6][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N0
cycloneive_lcell_comb \Mux9~11 (
// Equation(s):
// \Mux9~11_combout  = (\Mux9~10_combout  & ((\regs[7][22]~q ) # ((!dcifimemload_22)))) # (!\Mux9~10_combout  & (((\regs[6][22]~q  & dcifimemload_22))))

	.dataa(\Mux9~10_combout ),
	.datab(\regs[7][22]~q ),
	.datac(\regs[6][22]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~11 .lut_mask = 16'hD8AA;
defparam \Mux9~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N11
dffeas \regs[13][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][22] .is_wysiwyg = "true";
defparam \regs[13][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N10
cycloneive_lcell_comb \Mux9~17 (
// Equation(s):
// \Mux9~17_combout  = (dcifimemload_21 & (((\regs[13][22]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][22]~q  & ((!dcifimemload_22))))

	.dataa(\regs[12][22]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[13][22]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~17 .lut_mask = 16'hCCE2;
defparam \Mux9~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N4
cycloneive_lcell_comb \Mux9~18 (
// Equation(s):
// \Mux9~18_combout  = (\Mux9~17_combout  & ((\regs[15][22]~q ) # ((!dcifimemload_22)))) # (!\Mux9~17_combout  & (((\regs[14][22]~q  & dcifimemload_22))))

	.dataa(\regs[15][22]~q ),
	.datab(\regs[14][22]~q ),
	.datac(\Mux9~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~18 .lut_mask = 16'hACF0;
defparam \Mux9~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y45_N14
cycloneive_lcell_comb \regs[3][22]~feeder (
// Equation(s):
// \regs[3][22]~feeder_combout  = \regs~24_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~24_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[3][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][22]~feeder .lut_mask = 16'hF0F0;
defparam \regs[3][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y45_N15
dffeas \regs[3][22] (
	.clk(CLK),
	.d(\regs[3][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][22] .is_wysiwyg = "true";
defparam \regs[3][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y45_N20
cycloneive_lcell_comb \Mux9~14 (
// Equation(s):
// \Mux9~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][22]~q ))) # (!dcifimemload_22 & (\regs[1][22]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[1][22]~q ),
	.datac(\regs[3][22]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~14 .lut_mask = 16'hA088;
defparam \Mux9~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N30
cycloneive_lcell_comb \Mux9~15 (
// Equation(s):
// \Mux9~15_combout  = (\Mux9~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \regs[2][22]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[2][22]~q ),
	.datad(\Mux9~14_combout ),
	.cin(gnd),
	.combout(\Mux9~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~15 .lut_mask = 16'hFF40;
defparam \Mux9~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N1
dffeas \regs[8][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~24_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][22] .is_wysiwyg = "true";
defparam \regs[8][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N0
cycloneive_lcell_comb \Mux9~12 (
// Equation(s):
// \Mux9~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\regs[10][22]~q )) # (!dcifimemload_22 & ((\regs[8][22]~q )))))

	.dataa(\regs[10][22]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[8][22]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~12 .lut_mask = 16'hEE30;
defparam \Mux9~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N26
cycloneive_lcell_comb \Mux9~13 (
// Equation(s):
// \Mux9~13_combout  = (dcifimemload_21 & ((\Mux9~12_combout  & ((\regs[11][22]~q ))) # (!\Mux9~12_combout  & (\regs[9][22]~q )))) # (!dcifimemload_21 & (((\Mux9~12_combout ))))

	.dataa(\regs[9][22]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[11][22]~q ),
	.datad(\Mux9~12_combout ),
	.cin(gnd),
	.combout(\Mux9~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~13 .lut_mask = 16'hF388;
defparam \Mux9~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N24
cycloneive_lcell_comb \Mux9~16 (
// Equation(s):
// \Mux9~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux9~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & (\Mux9~15_combout )))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux9~15_combout ),
	.datad(\Mux9~13_combout ),
	.cin(gnd),
	.combout(\Mux9~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~16 .lut_mask = 16'hBA98;
defparam \Mux9~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N10
cycloneive_lcell_comb \Mux9~19 (
// Equation(s):
// \Mux9~19_combout  = (dcifimemload_23 & ((\Mux9~16_combout  & ((\Mux9~18_combout ))) # (!\Mux9~16_combout  & (\Mux9~11_combout )))) # (!dcifimemload_23 & (((\Mux9~16_combout ))))

	.dataa(\Mux9~11_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux9~18_combout ),
	.datad(\Mux9~16_combout ),
	.cin(gnd),
	.combout(\Mux9~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~19 .lut_mask = 16'hF388;
defparam \Mux9~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N18
cycloneive_lcell_comb \regs~25 (
// Equation(s):
// \regs~25_combout  = (\Selector10~1_combout  & !\Equal0~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector10),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\regs~25_combout ),
	.cout());
// synopsys translate_off
defparam \regs~25 .lut_mask = 16'h00F0;
defparam \regs~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N26
cycloneive_lcell_comb \regs[23][21]~feeder (
// Equation(s):
// \regs[23][21]~feeder_combout  = \regs~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~25_combout ),
	.cin(gnd),
	.combout(\regs[23][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][21]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N27
dffeas \regs[23][21] (
	.clk(CLK),
	.d(\regs[23][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][21] .is_wysiwyg = "true";
defparam \regs[23][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N7
dffeas \regs[31][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][21] .is_wysiwyg = "true";
defparam \regs[31][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N24
cycloneive_lcell_comb \regs[27][21]~feeder (
// Equation(s):
// \regs[27][21]~feeder_combout  = \regs~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~25_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][21]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N25
dffeas \regs[27][21] (
	.clk(CLK),
	.d(\regs[27][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][21] .is_wysiwyg = "true";
defparam \regs[27][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N10
cycloneive_lcell_comb \Mux42~7 (
// Equation(s):
// \Mux42~7_combout  = (dcifimemload_19 & (((\regs[27][21]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\regs[19][21]~q  & ((!dcifimemload_18))))

	.dataa(\regs[19][21]~q ),
	.datab(\regs[27][21]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux42~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~7 .lut_mask = 16'hF0CA;
defparam \Mux42~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N24
cycloneive_lcell_comb \Mux42~8 (
// Equation(s):
// \Mux42~8_combout  = (dcifimemload_18 & ((\Mux42~7_combout  & ((\regs[31][21]~q ))) # (!\Mux42~7_combout  & (\regs[23][21]~q )))) # (!dcifimemload_18 & (((\Mux42~7_combout ))))

	.dataa(\regs[23][21]~q ),
	.datab(\regs[31][21]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux42~7_combout ),
	.cin(gnd),
	.combout(\Mux42~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~8 .lut_mask = 16'hCFA0;
defparam \Mux42~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N10
cycloneive_lcell_comb \regs[21][21]~feeder (
// Equation(s):
// \regs[21][21]~feeder_combout  = \regs~25_combout 

	.dataa(gnd),
	.datab(\regs~25_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[21][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][21]~feeder .lut_mask = 16'hCCCC;
defparam \regs[21][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N11
dffeas \regs[21][21] (
	.clk(CLK),
	.d(\regs[21][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][21] .is_wysiwyg = "true";
defparam \regs[21][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N26
cycloneive_lcell_comb \regs[29][21]~feeder (
// Equation(s):
// \regs[29][21]~feeder_combout  = \regs~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~25_combout ),
	.cin(gnd),
	.combout(\regs[29][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][21]~feeder .lut_mask = 16'hFF00;
defparam \regs[29][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N27
dffeas \regs[29][21] (
	.clk(CLK),
	.d(\regs[29][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][21] .is_wysiwyg = "true";
defparam \regs[29][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N24
cycloneive_lcell_comb \regs[17][21]~feeder (
// Equation(s):
// \regs[17][21]~feeder_combout  = \regs~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~25_combout ),
	.cin(gnd),
	.combout(\regs[17][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][21]~feeder .lut_mask = 16'hFF00;
defparam \regs[17][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N25
dffeas \regs[17][21] (
	.clk(CLK),
	.d(\regs[17][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][21] .is_wysiwyg = "true";
defparam \regs[17][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N10
cycloneive_lcell_comb \regs[25][21]~feeder (
// Equation(s):
// \regs[25][21]~feeder_combout  = \regs~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~25_combout ),
	.cin(gnd),
	.combout(\regs[25][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[25][21]~feeder .lut_mask = 16'hFF00;
defparam \regs[25][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N11
dffeas \regs[25][21] (
	.clk(CLK),
	.d(\regs[25][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][21] .is_wysiwyg = "true";
defparam \regs[25][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N24
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[25][21]~q ))) # (!dcifimemload_19 & (\regs[17][21]~q ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\regs[17][21]~q ),
	.datad(\regs[25][21]~q ),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hDC98;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N4
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (\Mux42~0_combout  & (((\regs[29][21]~q ) # (!dcifimemload_18)))) # (!\Mux42~0_combout  & (\regs[21][21]~q  & ((dcifimemload_18))))

	.dataa(\regs[21][21]~q ),
	.datab(\regs[29][21]~q ),
	.datac(\Mux42~0_combout ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hCAF0;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N9
dffeas \regs[24][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][21] .is_wysiwyg = "true";
defparam \regs[24][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N3
dffeas \regs[20][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][21] .is_wysiwyg = "true";
defparam \regs[20][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N2
cycloneive_lcell_comb \Mux42~4 (
// Equation(s):
// \Mux42~4_combout  = (dcifimemload_18 & (((\regs[20][21]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[16][21]~q  & ((!dcifimemload_19))))

	.dataa(\regs[16][21]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[20][21]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux42~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~4 .lut_mask = 16'hCCE2;
defparam \Mux42~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N8
cycloneive_lcell_comb \Mux42~5 (
// Equation(s):
// \Mux42~5_combout  = (dcifimemload_19 & ((\Mux42~4_combout  & (\regs[28][21]~q )) # (!\Mux42~4_combout  & ((\regs[24][21]~q ))))) # (!dcifimemload_19 & (((\Mux42~4_combout ))))

	.dataa(\regs[28][21]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[24][21]~q ),
	.datad(\Mux42~4_combout ),
	.cin(gnd),
	.combout(\Mux42~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~5 .lut_mask = 16'hBBC0;
defparam \Mux42~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y43_N7
dffeas \regs[26][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][21] .is_wysiwyg = "true";
defparam \regs[26][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y43_N1
dffeas \regs[22][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][21] .is_wysiwyg = "true";
defparam \regs[22][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N0
cycloneive_lcell_comb \Mux42~2 (
// Equation(s):
// \Mux42~2_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\regs[22][21]~q ))) # (!dcifimemload_18 & (\regs[18][21]~q ))))

	.dataa(\regs[18][21]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[22][21]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux42~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~2 .lut_mask = 16'hFC22;
defparam \Mux42~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y43_N6
cycloneive_lcell_comb \Mux42~3 (
// Equation(s):
// \Mux42~3_combout  = (dcifimemload_19 & ((\Mux42~2_combout  & (\regs[30][21]~q )) # (!\Mux42~2_combout  & ((\regs[26][21]~q ))))) # (!dcifimemload_19 & (((\Mux42~2_combout ))))

	.dataa(\regs[30][21]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[26][21]~q ),
	.datad(\Mux42~2_combout ),
	.cin(gnd),
	.combout(\Mux42~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~3 .lut_mask = 16'hBBC0;
defparam \Mux42~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N6
cycloneive_lcell_comb \Mux42~6 (
// Equation(s):
// \Mux42~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux42~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux42~5_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux42~5_combout ),
	.datad(\Mux42~3_combout ),
	.cin(gnd),
	.combout(\Mux42~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~6 .lut_mask = 16'hBA98;
defparam \Mux42~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N2
cycloneive_lcell_comb \regs[3][21]~feeder (
// Equation(s):
// \regs[3][21]~feeder_combout  = \regs~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~25_combout ),
	.cin(gnd),
	.combout(\regs[3][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][21]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N3
dffeas \regs[3][21] (
	.clk(CLK),
	.d(\regs[3][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][21] .is_wysiwyg = "true";
defparam \regs[3][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y45_N5
dffeas \regs[1][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][21] .is_wysiwyg = "true";
defparam \regs[1][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N4
cycloneive_lcell_comb \Mux42~14 (
// Equation(s):
// \Mux42~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][21]~q )) # (!dcifimemload_17 & ((\regs[1][21]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[3][21]~q ),
	.datac(\regs[1][21]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux42~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~14 .lut_mask = 16'h88A0;
defparam \Mux42~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y45_N11
dffeas \regs[2][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][21] .is_wysiwyg = "true";
defparam \regs[2][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N10
cycloneive_lcell_comb \Mux42~15 (
// Equation(s):
// \Mux42~15_combout  = (\Mux42~14_combout ) # ((!dcifimemload_16 & (\regs[2][21]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\Mux42~14_combout ),
	.datac(\regs[2][21]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux42~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~15 .lut_mask = 16'hDCCC;
defparam \Mux42~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N24
cycloneive_lcell_comb \regs[9][21]~feeder (
// Equation(s):
// \regs[9][21]~feeder_combout  = \regs~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~25_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][21]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N25
dffeas \regs[9][21] (
	.clk(CLK),
	.d(\regs[9][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][21] .is_wysiwyg = "true";
defparam \regs[9][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N1
dffeas \regs[11][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][21] .is_wysiwyg = "true";
defparam \regs[11][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N4
cycloneive_lcell_comb \regs[8][21]~feeder (
// Equation(s):
// \regs[8][21]~feeder_combout  = \regs~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~25_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[8][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][21]~feeder .lut_mask = 16'hF0F0;
defparam \regs[8][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y32_N5
dffeas \regs[8][21] (
	.clk(CLK),
	.d(\regs[8][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][21] .is_wysiwyg = "true";
defparam \regs[8][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N18
cycloneive_lcell_comb \Mux42~12 (
// Equation(s):
// \Mux42~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][21]~q )) # (!dcifimemload_17 & ((\regs[8][21]~q )))))

	.dataa(\regs[10][21]~q ),
	.datab(\regs[8][21]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux42~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~12 .lut_mask = 16'hFA0C;
defparam \Mux42~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N0
cycloneive_lcell_comb \Mux42~13 (
// Equation(s):
// \Mux42~13_combout  = (dcifimemload_16 & ((\Mux42~12_combout  & ((\regs[11][21]~q ))) # (!\Mux42~12_combout  & (\regs[9][21]~q )))) # (!dcifimemload_16 & (((\Mux42~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][21]~q ),
	.datac(\regs[11][21]~q ),
	.datad(\Mux42~12_combout ),
	.cin(gnd),
	.combout(\Mux42~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~13 .lut_mask = 16'hF588;
defparam \Mux42~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N30
cycloneive_lcell_comb \Mux42~16 (
// Equation(s):
// \Mux42~16_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux42~13_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & (\Mux42~15_combout )))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux42~15_combout ),
	.datad(\Mux42~13_combout ),
	.cin(gnd),
	.combout(\Mux42~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~16 .lut_mask = 16'hBA98;
defparam \Mux42~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N31
dffeas \regs[5][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][21] .is_wysiwyg = "true";
defparam \regs[5][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N30
cycloneive_lcell_comb \Mux42~10 (
// Equation(s):
// \Mux42~10_combout  = (dcifimemload_16 & (((\regs[5][21]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][21]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][21]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[5][21]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux42~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~10 .lut_mask = 16'hCCE2;
defparam \Mux42~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N27
dffeas \regs[7][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][21] .is_wysiwyg = "true";
defparam \regs[7][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N1
dffeas \regs[6][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][21] .is_wysiwyg = "true";
defparam \regs[6][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N0
cycloneive_lcell_comb \Mux42~11 (
// Equation(s):
// \Mux42~11_combout  = (\Mux42~10_combout  & ((\regs[7][21]~q ) # ((!dcifimemload_17)))) # (!\Mux42~10_combout  & (((\regs[6][21]~q  & dcifimemload_17))))

	.dataa(\Mux42~10_combout ),
	.datab(\regs[7][21]~q ),
	.datac(\regs[6][21]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux42~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~11 .lut_mask = 16'hD8AA;
defparam \Mux42~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y44_N31
dffeas \regs[12][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][21] .is_wysiwyg = "true";
defparam \regs[12][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N30
cycloneive_lcell_comb \Mux42~17 (
// Equation(s):
// \Mux42~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][21]~q )) # (!dcifimemload_16 & ((\regs[12][21]~q )))))

	.dataa(\regs[13][21]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][21]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux42~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~17 .lut_mask = 16'hEE30;
defparam \Mux42~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y44_N1
dffeas \regs[14][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][21] .is_wysiwyg = "true";
defparam \regs[14][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y44_N15
dffeas \regs[15][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][21] .is_wysiwyg = "true";
defparam \regs[15][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N14
cycloneive_lcell_comb \Mux42~18 (
// Equation(s):
// \Mux42~18_combout  = (\Mux42~17_combout  & (((\regs[15][21]~q ) # (!dcifimemload_17)))) # (!\Mux42~17_combout  & (\regs[14][21]~q  & ((dcifimemload_17))))

	.dataa(\Mux42~17_combout ),
	.datab(\regs[14][21]~q ),
	.datac(\regs[15][21]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux42~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~18 .lut_mask = 16'hE4AA;
defparam \Mux42~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N16
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[21][21]~q ))) # (!dcifimemload_23 & (\regs[17][21]~q ))))

	.dataa(\regs[17][21]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[21][21]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hFC22;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N14
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (dcifimemload_24 & ((\Mux10~0_combout  & (\regs[29][21]~q )) # (!\Mux10~0_combout  & ((\regs[25][21]~q ))))) # (!dcifimemload_24 & (((\Mux10~0_combout ))))

	.dataa(\regs[29][21]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[25][21]~q ),
	.datad(\Mux10~0_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hBBC0;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N5
dffeas \regs[28][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][21] .is_wysiwyg = "true";
defparam \regs[28][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y42_N3
dffeas \regs[16][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][21] .is_wysiwyg = "true";
defparam \regs[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N2
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[24][21]~q )) # (!dcifimemload_24 & ((\regs[16][21]~q )))))

	.dataa(dcifimemload_23),
	.datab(\regs[24][21]~q ),
	.datac(\regs[16][21]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hEE50;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N4
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// \Mux10~5_combout  = (dcifimemload_23 & ((\Mux10~4_combout  & ((\regs[28][21]~q ))) # (!\Mux10~4_combout  & (\regs[20][21]~q )))) # (!dcifimemload_23 & (((\Mux10~4_combout ))))

	.dataa(\regs[20][21]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[28][21]~q ),
	.datad(\Mux10~4_combout ),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hF388;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N19
dffeas \regs[30][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][21] .is_wysiwyg = "true";
defparam \regs[30][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N18
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (\Mux10~2_combout  & (((\regs[30][21]~q ) # (!dcifimemload_23)))) # (!\Mux10~2_combout  & (\regs[22][21]~q  & ((dcifimemload_23))))

	.dataa(\Mux10~2_combout ),
	.datab(\regs[22][21]~q ),
	.datac(\regs[30][21]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hE4AA;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N8
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux10~3_combout ))) # (!dcifimemload_22 & (\Mux10~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux10~5_combout ),
	.datad(\Mux10~3_combout ),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hDC98;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N25
dffeas \regs[19][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][21] .is_wysiwyg = "true";
defparam \regs[19][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N24
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// \Mux10~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[23][21]~q )) # (!dcifimemload_23 & ((\regs[19][21]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[23][21]~q ),
	.datac(\regs[19][21]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hEE50;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N6
cycloneive_lcell_comb \Mux10~8 (
// Equation(s):
// \Mux10~8_combout  = (dcifimemload_24 & ((\Mux10~7_combout  & ((\regs[31][21]~q ))) # (!\Mux10~7_combout  & (\regs[27][21]~q )))) # (!dcifimemload_24 & (((\Mux10~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][21]~q ),
	.datac(\regs[31][21]~q ),
	.datad(\Mux10~7_combout ),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~8 .lut_mask = 16'hF588;
defparam \Mux10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N30
cycloneive_lcell_comb \Mux10~9 (
// Equation(s):
// \Mux10~9_combout  = (dcifimemload_21 & ((\Mux10~6_combout  & ((\Mux10~8_combout ))) # (!\Mux10~6_combout  & (\Mux10~1_combout )))) # (!dcifimemload_21 & (((\Mux10~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux10~1_combout ),
	.datac(\Mux10~6_combout ),
	.datad(\Mux10~8_combout ),
	.cin(gnd),
	.combout(\Mux10~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~9 .lut_mask = 16'hF858;
defparam \Mux10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y44_N29
dffeas \regs[13][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][21] .is_wysiwyg = "true";
defparam \regs[13][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N28
cycloneive_lcell_comb \Mux10~17 (
// Equation(s):
// \Mux10~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\regs[13][21]~q ))) # (!dcifimemload_21 & (\regs[12][21]~q ))))

	.dataa(\regs[12][21]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[13][21]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux10~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~17 .lut_mask = 16'hFC22;
defparam \Mux10~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N0
cycloneive_lcell_comb \Mux10~18 (
// Equation(s):
// \Mux10~18_combout  = (dcifimemload_22 & ((\Mux10~17_combout  & (\regs[15][21]~q )) # (!\Mux10~17_combout  & ((\regs[14][21]~q ))))) # (!dcifimemload_22 & (((\Mux10~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][21]~q ),
	.datac(\regs[14][21]~q ),
	.datad(\Mux10~17_combout ),
	.cin(gnd),
	.combout(\Mux10~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~18 .lut_mask = 16'hDDA0;
defparam \Mux10~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N23
dffeas \regs[10][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][21] .is_wysiwyg = "true";
defparam \regs[10][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \Mux10~10 (
// Equation(s):
// \Mux10~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][21]~q ))) # (!dcifimemload_22 & (\regs[8][21]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][21]~q ),
	.datac(\regs[10][21]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux10~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~10 .lut_mask = 16'hFA44;
defparam \Mux10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N2
cycloneive_lcell_comb \Mux10~11 (
// Equation(s):
// \Mux10~11_combout  = (\Mux10~10_combout  & ((\regs[11][21]~q ) # ((!dcifimemload_21)))) # (!\Mux10~10_combout  & (((\regs[9][21]~q  & dcifimemload_21))))

	.dataa(\regs[11][21]~q ),
	.datab(\regs[9][21]~q ),
	.datac(\Mux10~10_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~11 .lut_mask = 16'hACF0;
defparam \Mux10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N16
cycloneive_lcell_comb \Mux10~14 (
// Equation(s):
// \Mux10~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\regs[3][21]~q )) # (!dcifimemload_22 & ((\regs[1][21]~q )))))

	.dataa(dcifimemload_21),
	.datab(\regs[3][21]~q ),
	.datac(\regs[1][21]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux10~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~14 .lut_mask = 16'h88A0;
defparam \Mux10~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N18
cycloneive_lcell_comb \Mux10~15 (
// Equation(s):
// \Mux10~15_combout  = (\Mux10~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \regs[2][21]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[2][21]~q ),
	.datad(\Mux10~14_combout ),
	.cin(gnd),
	.combout(\Mux10~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~15 .lut_mask = 16'hFF40;
defparam \Mux10~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N29
dffeas \regs[4][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][21] .is_wysiwyg = "true";
defparam \regs[4][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N28
cycloneive_lcell_comb \Mux10~12 (
// Equation(s):
// \Mux10~12_combout  = (dcifimemload_21 & ((dcifimemload_22) # ((\regs[5][21]~q )))) # (!dcifimemload_21 & (!dcifimemload_22 & (\regs[4][21]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[4][21]~q ),
	.datad(\regs[5][21]~q ),
	.cin(gnd),
	.combout(\Mux10~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~12 .lut_mask = 16'hBA98;
defparam \Mux10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N26
cycloneive_lcell_comb \Mux10~13 (
// Equation(s):
// \Mux10~13_combout  = (dcifimemload_22 & ((\Mux10~12_combout  & ((\regs[7][21]~q ))) # (!\Mux10~12_combout  & (\regs[6][21]~q )))) # (!dcifimemload_22 & (((\Mux10~12_combout ))))

	.dataa(\regs[6][21]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[7][21]~q ),
	.datad(\Mux10~12_combout ),
	.cin(gnd),
	.combout(\Mux10~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~13 .lut_mask = 16'hF388;
defparam \Mux10~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N24
cycloneive_lcell_comb \Mux10~16 (
// Equation(s):
// \Mux10~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux10~13_combout ))) # (!dcifimemload_23 & (\Mux10~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux10~15_combout ),
	.datad(\Mux10~13_combout ),
	.cin(gnd),
	.combout(\Mux10~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~16 .lut_mask = 16'hDC98;
defparam \Mux10~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N18
cycloneive_lcell_comb \Mux10~19 (
// Equation(s):
// \Mux10~19_combout  = (dcifimemload_24 & ((\Mux10~16_combout  & (\Mux10~18_combout )) # (!\Mux10~16_combout  & ((\Mux10~11_combout ))))) # (!dcifimemload_24 & (((\Mux10~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux10~18_combout ),
	.datac(\Mux10~11_combout ),
	.datad(\Mux10~16_combout ),
	.cin(gnd),
	.combout(\Mux10~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~19 .lut_mask = 16'hDDA0;
defparam \Mux10~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N24
cycloneive_lcell_comb \regs~26 (
// Equation(s):
// \regs~26_combout  = (!\Equal0~1_combout  & \Selector11~1_combout )

	.dataa(\Equal0~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector11),
	.cin(gnd),
	.combout(\regs~26_combout ),
	.cout());
// synopsys translate_off
defparam \regs~26 .lut_mask = 16'h5500;
defparam \regs~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N28
cycloneive_lcell_comb \regs[27][20]~feeder (
// Equation(s):
// \regs[27][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~26_combout ),
	.cin(gnd),
	.combout(\regs[27][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][20]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y45_N29
dffeas \regs[27][20] (
	.clk(CLK),
	.d(\regs[27][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][20] .is_wysiwyg = "true";
defparam \regs[27][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N17
dffeas \regs[31][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][20] .is_wysiwyg = "true";
defparam \regs[31][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N11
dffeas \regs[23][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][20] .is_wysiwyg = "true";
defparam \regs[23][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N19
dffeas \regs[19][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][20] .is_wysiwyg = "true";
defparam \regs[19][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N18
cycloneive_lcell_comb \Mux43~7 (
// Equation(s):
// \Mux43~7_combout  = (dcifimemload_18 & ((\regs[23][20]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[19][20]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[23][20]~q ),
	.datac(\regs[19][20]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux43~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~7 .lut_mask = 16'hAAD8;
defparam \Mux43~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N16
cycloneive_lcell_comb \Mux43~8 (
// Equation(s):
// \Mux43~8_combout  = (dcifimemload_19 & ((\Mux43~7_combout  & ((\regs[31][20]~q ))) # (!\Mux43~7_combout  & (\regs[27][20]~q )))) # (!dcifimemload_19 & (((\Mux43~7_combout ))))

	.dataa(\regs[27][20]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[31][20]~q ),
	.datad(\Mux43~7_combout ),
	.cin(gnd),
	.combout(\Mux43~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~8 .lut_mask = 16'hF388;
defparam \Mux43~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N31
dffeas \regs[28][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][20] .is_wysiwyg = "true";
defparam \regs[28][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N17
dffeas \regs[16][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][20] .is_wysiwyg = "true";
defparam \regs[16][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N16
cycloneive_lcell_comb \Mux43~4 (
// Equation(s):
// \Mux43~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[24][20]~q )) # (!dcifimemload_19 & ((\regs[16][20]~q )))))

	.dataa(\regs[24][20]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[16][20]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux43~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~4 .lut_mask = 16'hEE30;
defparam \Mux43~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N30
cycloneive_lcell_comb \Mux43~5 (
// Equation(s):
// \Mux43~5_combout  = (dcifimemload_18 & ((\Mux43~4_combout  & ((\regs[28][20]~q ))) # (!\Mux43~4_combout  & (\regs[20][20]~q )))) # (!dcifimemload_18 & (((\Mux43~4_combout ))))

	.dataa(\regs[20][20]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[28][20]~q ),
	.datad(\Mux43~4_combout ),
	.cin(gnd),
	.combout(\Mux43~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~5 .lut_mask = 16'hF388;
defparam \Mux43~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N17
dffeas \regs[30][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][20] .is_wysiwyg = "true";
defparam \regs[30][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N19
dffeas \regs[18][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][20] .is_wysiwyg = "true";
defparam \regs[18][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N18
cycloneive_lcell_comb \Mux43~2 (
// Equation(s):
// \Mux43~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[26][20]~q )) # (!dcifimemload_19 & ((\regs[18][20]~q )))))

	.dataa(\regs[26][20]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][20]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux43~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~2 .lut_mask = 16'hEE30;
defparam \Mux43~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N16
cycloneive_lcell_comb \Mux43~3 (
// Equation(s):
// \Mux43~3_combout  = (dcifimemload_18 & ((\Mux43~2_combout  & ((\regs[30][20]~q ))) # (!\Mux43~2_combout  & (\regs[22][20]~q )))) # (!dcifimemload_18 & (((\Mux43~2_combout ))))

	.dataa(\regs[22][20]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[30][20]~q ),
	.datad(\Mux43~2_combout ),
	.cin(gnd),
	.combout(\Mux43~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~3 .lut_mask = 16'hF388;
defparam \Mux43~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N4
cycloneive_lcell_comb \Mux43~6 (
// Equation(s):
// \Mux43~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux43~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux43~5_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux43~5_combout ),
	.datad(\Mux43~3_combout ),
	.cin(gnd),
	.combout(\Mux43~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~6 .lut_mask = 16'hBA98;
defparam \Mux43~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N25
dffeas \regs[25][20] (
	.clk(CLK),
	.d(\regs~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][20] .is_wysiwyg = "true";
defparam \regs[25][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N6
cycloneive_lcell_comb \regs[29][20]~feeder (
// Equation(s):
// \regs[29][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~26_combout ),
	.cin(gnd),
	.combout(\regs[29][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][20]~feeder .lut_mask = 16'hFF00;
defparam \regs[29][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N7
dffeas \regs[29][20] (
	.clk(CLK),
	.d(\regs[29][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][20] .is_wysiwyg = "true";
defparam \regs[29][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N0
cycloneive_lcell_comb \regs[21][20]~feeder (
// Equation(s):
// \regs[21][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~26_combout ),
	.cin(gnd),
	.combout(\regs[21][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][20]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N1
dffeas \regs[21][20] (
	.clk(CLK),
	.d(\regs[21][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][20] .is_wysiwyg = "true";
defparam \regs[21][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N13
dffeas \regs[17][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][20] .is_wysiwyg = "true";
defparam \regs[17][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N12
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[21][20]~q )) # (!dcifimemload_18 & ((\regs[17][20]~q )))))

	.dataa(dcifimemload_19),
	.datab(\regs[21][20]~q ),
	.datac(\regs[17][20]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hEE50;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N28
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (dcifimemload_19 & ((\Mux43~0_combout  & ((\regs[29][20]~q ))) # (!\Mux43~0_combout  & (\regs[25][20]~q )))) # (!dcifimemload_19 & (((\Mux43~0_combout ))))

	.dataa(\regs[25][20]~q ),
	.datab(\regs[29][20]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux43~0_combout ),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hCFA0;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N20
cycloneive_lcell_comb \regs[14][20]~feeder (
// Equation(s):
// \regs[14][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~26_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[14][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][20]~feeder .lut_mask = 16'hF0F0;
defparam \regs[14][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y44_N21
dffeas \regs[14][20] (
	.clk(CLK),
	.d(\regs[14][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][20] .is_wysiwyg = "true";
defparam \regs[14][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y44_N7
dffeas \regs[15][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][20] .is_wysiwyg = "true";
defparam \regs[15][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y44_N7
dffeas \regs[12][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][20] .is_wysiwyg = "true";
defparam \regs[12][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N6
cycloneive_lcell_comb \Mux43~17 (
// Equation(s):
// \Mux43~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][20]~q )) # (!dcifimemload_16 & ((\regs[12][20]~q )))))

	.dataa(\regs[13][20]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][20]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux43~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~17 .lut_mask = 16'hEE30;
defparam \Mux43~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N6
cycloneive_lcell_comb \Mux43~18 (
// Equation(s):
// \Mux43~18_combout  = (dcifimemload_17 & ((\Mux43~17_combout  & ((\regs[15][20]~q ))) # (!\Mux43~17_combout  & (\regs[14][20]~q )))) # (!dcifimemload_17 & (((\Mux43~17_combout ))))

	.dataa(\regs[14][20]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[15][20]~q ),
	.datad(\Mux43~17_combout ),
	.cin(gnd),
	.combout(\Mux43~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~18 .lut_mask = 16'hF388;
defparam \Mux43~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N30
cycloneive_lcell_comb \regs[9][20]~feeder (
// Equation(s):
// \regs[9][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~26_combout ),
	.cin(gnd),
	.combout(\regs[9][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][20]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N31
dffeas \regs[9][20] (
	.clk(CLK),
	.d(\regs[9][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][20] .is_wysiwyg = "true";
defparam \regs[9][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N9
dffeas \regs[11][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][20] .is_wysiwyg = "true";
defparam \regs[11][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \regs[8][20]~feeder (
// Equation(s):
// \regs[8][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~26_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[8][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][20]~feeder .lut_mask = 16'hF0F0;
defparam \regs[8][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N3
dffeas \regs[8][20] (
	.clk(CLK),
	.d(\regs[8][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][20] .is_wysiwyg = "true";
defparam \regs[8][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N29
dffeas \regs[10][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][20] .is_wysiwyg = "true";
defparam \regs[10][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N18
cycloneive_lcell_comb \Mux43~10 (
// Equation(s):
// \Mux43~10_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\regs[10][20]~q ))) # (!dcifimemload_17 & (\regs[8][20]~q ))))

	.dataa(dcifimemload_16),
	.datab(\regs[8][20]~q ),
	.datac(\regs[10][20]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux43~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~10 .lut_mask = 16'hFA44;
defparam \Mux43~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N8
cycloneive_lcell_comb \Mux43~11 (
// Equation(s):
// \Mux43~11_combout  = (dcifimemload_16 & ((\Mux43~10_combout  & ((\regs[11][20]~q ))) # (!\Mux43~10_combout  & (\regs[9][20]~q )))) # (!dcifimemload_16 & (((\Mux43~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][20]~q ),
	.datac(\regs[11][20]~q ),
	.datad(\Mux43~10_combout ),
	.cin(gnd),
	.combout(\Mux43~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~11 .lut_mask = 16'hF588;
defparam \Mux43~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y45_N31
dffeas \regs[2][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][20] .is_wysiwyg = "true";
defparam \regs[2][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y45_N13
dffeas \regs[1][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][20] .is_wysiwyg = "true";
defparam \regs[1][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N12
cycloneive_lcell_comb \Mux43~14 (
// Equation(s):
// \Mux43~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][20]~q )) # (!dcifimemload_17 & ((\regs[1][20]~q )))))

	.dataa(\regs[3][20]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][20]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux43~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~14 .lut_mask = 16'h88C0;
defparam \Mux43~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N30
cycloneive_lcell_comb \Mux43~15 (
// Equation(s):
// \Mux43~15_combout  = (\Mux43~14_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][20]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[2][20]~q ),
	.datad(\Mux43~14_combout ),
	.cin(gnd),
	.combout(\Mux43~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~15 .lut_mask = 16'hFF20;
defparam \Mux43~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y45_N28
cycloneive_lcell_comb \regs[6][20]~feeder (
// Equation(s):
// \regs[6][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~26_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[6][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][20]~feeder .lut_mask = 16'hF0F0;
defparam \regs[6][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y45_N29
dffeas \regs[6][20] (
	.clk(CLK),
	.d(\regs[6][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][20] .is_wysiwyg = "true";
defparam \regs[6][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N11
dffeas \regs[7][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][20] .is_wysiwyg = "true";
defparam \regs[7][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N4
cycloneive_lcell_comb \regs[5][20]~feeder (
// Equation(s):
// \regs[5][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~26_combout ),
	.cin(gnd),
	.combout(\regs[5][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][20]~feeder .lut_mask = 16'hFF00;
defparam \regs[5][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N5
dffeas \regs[5][20] (
	.clk(CLK),
	.d(\regs[5][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][20] .is_wysiwyg = "true";
defparam \regs[5][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N17
dffeas \regs[4][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][20] .is_wysiwyg = "true";
defparam \regs[4][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N16
cycloneive_lcell_comb \Mux43~12 (
// Equation(s):
// \Mux43~12_combout  = (dcifimemload_16 & ((\regs[5][20]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][20]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[5][20]~q ),
	.datac(\regs[4][20]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux43~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~12 .lut_mask = 16'hAAD8;
defparam \Mux43~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N10
cycloneive_lcell_comb \Mux43~13 (
// Equation(s):
// \Mux43~13_combout  = (dcifimemload_17 & ((\Mux43~12_combout  & ((\regs[7][20]~q ))) # (!\Mux43~12_combout  & (\regs[6][20]~q )))) # (!dcifimemload_17 & (((\Mux43~12_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][20]~q ),
	.datac(\regs[7][20]~q ),
	.datad(\Mux43~12_combout ),
	.cin(gnd),
	.combout(\Mux43~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~13 .lut_mask = 16'hF588;
defparam \Mux43~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N24
cycloneive_lcell_comb \Mux43~16 (
// Equation(s):
// \Mux43~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux43~13_combout ))) # (!dcifimemload_18 & (\Mux43~15_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux43~15_combout ),
	.datad(\Mux43~13_combout ),
	.cin(gnd),
	.combout(\Mux43~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~16 .lut_mask = 16'hDC98;
defparam \Mux43~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N18
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// \Mux11~7_combout  = (dcifimemload_24 & (((\regs[27][20]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[19][20]~q  & ((!dcifimemload_23))))

	.dataa(\regs[19][20]~q ),
	.datab(\regs[27][20]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hF0CA;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N20
cycloneive_lcell_comb \Mux11~8 (
// Equation(s):
// \Mux11~8_combout  = (dcifimemload_23 & ((\Mux11~7_combout  & ((\regs[31][20]~q ))) # (!\Mux11~7_combout  & (\regs[23][20]~q )))) # (!dcifimemload_23 & (((\Mux11~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[23][20]~q ),
	.datac(\regs[31][20]~q ),
	.datad(\Mux11~7_combout ),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~8 .lut_mask = 16'hF588;
defparam \Mux11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N8
cycloneive_lcell_comb \regs[24][20]~feeder (
// Equation(s):
// \regs[24][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~26_combout ),
	.cin(gnd),
	.combout(\regs[24][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][20]~feeder .lut_mask = 16'hFF00;
defparam \regs[24][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N9
dffeas \regs[24][20] (
	.clk(CLK),
	.d(\regs[24][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][20] .is_wysiwyg = "true";
defparam \regs[24][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N9
dffeas \regs[20][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][20] .is_wysiwyg = "true";
defparam \regs[20][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N8
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[20][20]~q ))) # (!dcifimemload_23 & (\regs[16][20]~q ))))

	.dataa(dcifimemload_24),
	.datab(\regs[16][20]~q ),
	.datac(\regs[20][20]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hFA44;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N2
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// \Mux11~5_combout  = (\Mux11~4_combout  & ((\regs[28][20]~q ) # ((!dcifimemload_24)))) # (!\Mux11~4_combout  & (((\regs[24][20]~q  & dcifimemload_24))))

	.dataa(\regs[28][20]~q ),
	.datab(\regs[24][20]~q ),
	.datac(\Mux11~4_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hACF0;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y45_N13
dffeas \regs[26][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][20] .is_wysiwyg = "true";
defparam \regs[26][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N17
dffeas \regs[22][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][20] .is_wysiwyg = "true";
defparam \regs[22][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N16
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (dcifimemload_23 & (((\regs[22][20]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[18][20]~q  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[18][20]~q ),
	.datac(\regs[22][20]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hAAE4;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y45_N12
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (dcifimemload_24 & ((\Mux11~2_combout  & (\regs[30][20]~q )) # (!\Mux11~2_combout  & ((\regs[26][20]~q ))))) # (!dcifimemload_24 & (((\Mux11~2_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[30][20]~q ),
	.datac(\regs[26][20]~q ),
	.datad(\Mux11~2_combout ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hDDA0;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N8
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux11~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux11~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux11~5_combout ),
	.datad(\Mux11~3_combout ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hBA98;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N2
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (dcifimemload_24 & ((\regs[25][20]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[17][20]~q  & !dcifimemload_23))))

	.dataa(\regs[25][20]~q ),
	.datab(\regs[17][20]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hF0AC;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N20
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (dcifimemload_23 & ((\Mux11~0_combout  & (\regs[29][20]~q )) # (!\Mux11~0_combout  & ((\regs[21][20]~q ))))) # (!dcifimemload_23 & (((\Mux11~0_combout ))))

	.dataa(\regs[29][20]~q ),
	.datab(\regs[21][20]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hAFC0;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N14
cycloneive_lcell_comb \Mux11~9 (
// Equation(s):
// \Mux11~9_combout  = (dcifimemload_21 & ((\Mux11~6_combout  & (\Mux11~8_combout )) # (!\Mux11~6_combout  & ((\Mux11~1_combout ))))) # (!dcifimemload_21 & (((\Mux11~6_combout ))))

	.dataa(\Mux11~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux11~6_combout ),
	.datad(\Mux11~1_combout ),
	.cin(gnd),
	.combout(\Mux11~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~9 .lut_mask = 16'hBCB0;
defparam \Mux11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y45_N22
cycloneive_lcell_comb \Mux11~10 (
// Equation(s):
// \Mux11~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\regs[5][20]~q )) # (!dcifimemload_21 & ((\regs[4][20]~q )))))

	.dataa(\regs[5][20]~q ),
	.datab(\regs[4][20]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~10 .lut_mask = 16'hFA0C;
defparam \Mux11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y45_N20
cycloneive_lcell_comb \Mux11~11 (
// Equation(s):
// \Mux11~11_combout  = (dcifimemload_22 & ((\Mux11~10_combout  & (\regs[7][20]~q )) # (!\Mux11~10_combout  & ((\regs[6][20]~q ))))) # (!dcifimemload_22 & (((\Mux11~10_combout ))))

	.dataa(\regs[7][20]~q ),
	.datab(\regs[6][20]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux11~10_combout ),
	.cin(gnd),
	.combout(\Mux11~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~11 .lut_mask = 16'hAFC0;
defparam \Mux11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N0
cycloneive_lcell_comb \regs[13][20]~feeder (
// Equation(s):
// \regs[13][20]~feeder_combout  = \regs~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~26_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[13][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][20]~feeder .lut_mask = 16'hF0F0;
defparam \regs[13][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y44_N1
dffeas \regs[13][20] (
	.clk(CLK),
	.d(\regs[13][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][20] .is_wysiwyg = "true";
defparam \regs[13][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N8
cycloneive_lcell_comb \Mux11~17 (
// Equation(s):
// \Mux11~17_combout  = (dcifimemload_21 & (((\regs[13][20]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][20]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][20]~q ),
	.datac(\regs[13][20]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux11~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~17 .lut_mask = 16'hAAE4;
defparam \Mux11~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N6
cycloneive_lcell_comb \Mux11~18 (
// Equation(s):
// \Mux11~18_combout  = (\Mux11~17_combout  & (((\regs[15][20]~q ) # (!dcifimemload_22)))) # (!\Mux11~17_combout  & (\regs[14][20]~q  & ((dcifimemload_22))))

	.dataa(\regs[14][20]~q ),
	.datab(\regs[15][20]~q ),
	.datac(\Mux11~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux11~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~18 .lut_mask = 16'hCAF0;
defparam \Mux11~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N3
dffeas \regs[3][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~26_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][20] .is_wysiwyg = "true";
defparam \regs[3][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N4
cycloneive_lcell_comb \Mux11~14 (
// Equation(s):
// \Mux11~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\regs[3][20]~q )) # (!dcifimemload_22 & ((\regs[1][20]~q )))))

	.dataa(dcifimemload_21),
	.datab(\regs[3][20]~q ),
	.datac(\regs[1][20]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux11~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~14 .lut_mask = 16'h88A0;
defparam \Mux11~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N24
cycloneive_lcell_comb \Mux11~15 (
// Equation(s):
// \Mux11~15_combout  = (\Mux11~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][20]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[2][20]~q ),
	.datad(\Mux11~14_combout ),
	.cin(gnd),
	.combout(\Mux11~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~15 .lut_mask = 16'hFF20;
defparam \Mux11~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \Mux11~12 (
// Equation(s):
// \Mux11~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][20]~q ))) # (!dcifimemload_22 & (\regs[8][20]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][20]~q ),
	.datac(\regs[10][20]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux11~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~12 .lut_mask = 16'hFA44;
defparam \Mux11~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N26
cycloneive_lcell_comb \Mux11~13 (
// Equation(s):
// \Mux11~13_combout  = (\Mux11~12_combout  & (((\regs[11][20]~q ) # (!dcifimemload_21)))) # (!\Mux11~12_combout  & (\regs[9][20]~q  & ((dcifimemload_21))))

	.dataa(\regs[9][20]~q ),
	.datab(\regs[11][20]~q ),
	.datac(\Mux11~12_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux11~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~13 .lut_mask = 16'hCAF0;
defparam \Mux11~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N2
cycloneive_lcell_comb \Mux11~16 (
// Equation(s):
// \Mux11~16_combout  = (dcifimemload_24 & (((dcifimemload_23) # (\Mux11~13_combout )))) # (!dcifimemload_24 & (\Mux11~15_combout  & (!dcifimemload_23)))

	.dataa(dcifimemload_24),
	.datab(\Mux11~15_combout ),
	.datac(dcifimemload_23),
	.datad(\Mux11~13_combout ),
	.cin(gnd),
	.combout(\Mux11~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~16 .lut_mask = 16'hAEA4;
defparam \Mux11~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N28
cycloneive_lcell_comb \Mux11~19 (
// Equation(s):
// \Mux11~19_combout  = (dcifimemload_23 & ((\Mux11~16_combout  & ((\Mux11~18_combout ))) # (!\Mux11~16_combout  & (\Mux11~11_combout )))) # (!dcifimemload_23 & (((\Mux11~16_combout ))))

	.dataa(\Mux11~11_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux11~18_combout ),
	.datad(\Mux11~16_combout ),
	.cin(gnd),
	.combout(\Mux11~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~19 .lut_mask = 16'hF388;
defparam \Mux11~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N14
cycloneive_lcell_comb \regs~27 (
// Equation(s):
// \regs~27_combout  = (!\Equal0~1_combout  & \Selector12~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Equal0~1_combout ),
	.datad(Selector12),
	.cin(gnd),
	.combout(\regs~27_combout ),
	.cout());
// synopsys translate_off
defparam \regs~27 .lut_mask = 16'h0F00;
defparam \regs~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N23
dffeas \regs[23][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][19] .is_wysiwyg = "true";
defparam \regs[23][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N15
dffeas \regs[31][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][19] .is_wysiwyg = "true";
defparam \regs[31][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N20
cycloneive_lcell_comb \regs[27][19]~feeder (
// Equation(s):
// \regs[27][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~27_combout ),
	.cin(gnd),
	.combout(\regs[27][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N21
dffeas \regs[27][19] (
	.clk(CLK),
	.d(\regs[27][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][19] .is_wysiwyg = "true";
defparam \regs[27][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N24
cycloneive_lcell_comb \Mux44~7 (
// Equation(s):
// \Mux44~7_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[27][19]~q ))) # (!dcifimemload_19 & (\regs[19][19]~q ))))

	.dataa(\regs[19][19]~q ),
	.datab(\regs[27][19]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux44~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~7 .lut_mask = 16'hFC0A;
defparam \Mux44~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N14
cycloneive_lcell_comb \Mux44~8 (
// Equation(s):
// \Mux44~8_combout  = (dcifimemload_18 & ((\Mux44~7_combout  & ((\regs[31][19]~q ))) # (!\Mux44~7_combout  & (\regs[23][19]~q )))) # (!dcifimemload_18 & (((\Mux44~7_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[23][19]~q ),
	.datac(\regs[31][19]~q ),
	.datad(\Mux44~7_combout ),
	.cin(gnd),
	.combout(\Mux44~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~8 .lut_mask = 16'hF588;
defparam \Mux44~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N26
cycloneive_lcell_comb \regs[24][19]~feeder (
// Equation(s):
// \regs[24][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~27_combout ),
	.cin(gnd),
	.combout(\regs[24][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[24][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N27
dffeas \regs[24][19] (
	.clk(CLK),
	.d(\regs[24][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][19] .is_wysiwyg = "true";
defparam \regs[24][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N31
dffeas \regs[28][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][19] .is_wysiwyg = "true";
defparam \regs[28][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N25
dffeas \regs[16][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][19] .is_wysiwyg = "true";
defparam \regs[16][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N24
cycloneive_lcell_comb \Mux44~4 (
// Equation(s):
// \Mux44~4_combout  = (dcifimemload_18 & ((\regs[20][19]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[16][19]~q  & !dcifimemload_19))))

	.dataa(\regs[20][19]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[16][19]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux44~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~4 .lut_mask = 16'hCCB8;
defparam \Mux44~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N30
cycloneive_lcell_comb \Mux44~5 (
// Equation(s):
// \Mux44~5_combout  = (dcifimemload_19 & ((\Mux44~4_combout  & ((\regs[28][19]~q ))) # (!\Mux44~4_combout  & (\regs[24][19]~q )))) # (!dcifimemload_19 & (((\Mux44~4_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[24][19]~q ),
	.datac(\regs[28][19]~q ),
	.datad(\Mux44~4_combout ),
	.cin(gnd),
	.combout(\Mux44~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~5 .lut_mask = 16'hF588;
defparam \Mux44~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N9
dffeas \regs[26][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][19] .is_wysiwyg = "true";
defparam \regs[26][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N19
dffeas \regs[30][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][19] .is_wysiwyg = "true";
defparam \regs[30][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N25
dffeas \regs[18][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][19] .is_wysiwyg = "true";
defparam \regs[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N24
cycloneive_lcell_comb \Mux44~2 (
// Equation(s):
// \Mux44~2_combout  = (dcifimemload_18 & ((\regs[22][19]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[18][19]~q  & !dcifimemload_19))))

	.dataa(\regs[22][19]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][19]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux44~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~2 .lut_mask = 16'hCCB8;
defparam \Mux44~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N18
cycloneive_lcell_comb \Mux44~3 (
// Equation(s):
// \Mux44~3_combout  = (dcifimemload_19 & ((\Mux44~2_combout  & ((\regs[30][19]~q ))) # (!\Mux44~2_combout  & (\regs[26][19]~q )))) # (!dcifimemload_19 & (((\Mux44~2_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[26][19]~q ),
	.datac(\regs[30][19]~q ),
	.datad(\Mux44~2_combout ),
	.cin(gnd),
	.combout(\Mux44~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~3 .lut_mask = 16'hF588;
defparam \Mux44~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N8
cycloneive_lcell_comb \Mux44~6 (
// Equation(s):
// \Mux44~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux44~3_combout ))) # (!dcifimemload_17 & (\Mux44~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux44~5_combout ),
	.datad(\Mux44~3_combout ),
	.cin(gnd),
	.combout(\Mux44~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~6 .lut_mask = 16'hDC98;
defparam \Mux44~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N12
cycloneive_lcell_comb \regs[29][19]~feeder (
// Equation(s):
// \regs[29][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~27_combout ),
	.cin(gnd),
	.combout(\regs[29][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[29][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N13
dffeas \regs[29][19] (
	.clk(CLK),
	.d(\regs[29][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][19] .is_wysiwyg = "true";
defparam \regs[29][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N5
dffeas \regs[21][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][19] .is_wysiwyg = "true";
defparam \regs[21][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N6
cycloneive_lcell_comb \regs[25][19]~feeder (
// Equation(s):
// \regs[25][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~27_combout ),
	.cin(gnd),
	.combout(\regs[25][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[25][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[25][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N7
dffeas \regs[25][19] (
	.clk(CLK),
	.d(\regs[25][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][19] .is_wysiwyg = "true";
defparam \regs[25][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N25
dffeas \regs[17][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][19] .is_wysiwyg = "true";
defparam \regs[17][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N24
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (dcifimemload_19 & ((\regs[25][19]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\regs[17][19]~q  & !dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\regs[25][19]~q ),
	.datac(\regs[17][19]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hAAD8;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N10
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (dcifimemload_18 & ((\Mux44~0_combout  & (\regs[29][19]~q )) # (!\Mux44~0_combout  & ((\regs[21][19]~q ))))) # (!dcifimemload_18 & (((\Mux44~0_combout ))))

	.dataa(\regs[29][19]~q ),
	.datab(\regs[21][19]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux44~0_combout ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hAFC0;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N1
dffeas \regs[14][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][19] .is_wysiwyg = "true";
defparam \regs[14][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N17
dffeas \regs[15][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][19] .is_wysiwyg = "true";
defparam \regs[15][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N19
dffeas \regs[13][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][19] .is_wysiwyg = "true";
defparam \regs[13][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N24
cycloneive_lcell_comb \Mux44~17 (
// Equation(s):
// \Mux44~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\regs[13][19]~q ))) # (!dcifimemload_16 & (\regs[12][19]~q ))))

	.dataa(\regs[12][19]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[13][19]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux44~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~17 .lut_mask = 16'hFC22;
defparam \Mux44~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N16
cycloneive_lcell_comb \Mux44~18 (
// Equation(s):
// \Mux44~18_combout  = (dcifimemload_17 & ((\Mux44~17_combout  & ((\regs[15][19]~q ))) # (!\Mux44~17_combout  & (\regs[14][19]~q )))) # (!dcifimemload_17 & (((\Mux44~17_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[14][19]~q ),
	.datac(\regs[15][19]~q ),
	.datad(\Mux44~17_combout ),
	.cin(gnd),
	.combout(\Mux44~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~18 .lut_mask = 16'hF588;
defparam \Mux44~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y32_N27
dffeas \regs[2][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][19] .is_wysiwyg = "true";
defparam \regs[2][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N17
dffeas \regs[3][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][19] .is_wysiwyg = "true";
defparam \regs[3][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N1
dffeas \regs[1][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][19] .is_wysiwyg = "true";
defparam \regs[1][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N0
cycloneive_lcell_comb \Mux44~14 (
// Equation(s):
// \Mux44~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][19]~q )) # (!dcifimemload_17 & ((\regs[1][19]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[3][19]~q ),
	.datac(\regs[1][19]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux44~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~14 .lut_mask = 16'h88A0;
defparam \Mux44~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N26
cycloneive_lcell_comb \Mux44~15 (
// Equation(s):
// \Mux44~15_combout  = (\Mux44~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][19]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][19]~q ),
	.datad(\Mux44~14_combout ),
	.cin(gnd),
	.combout(\Mux44~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~15 .lut_mask = 16'hFF40;
defparam \Mux44~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N8
cycloneive_lcell_comb \regs[9][19]~feeder (
// Equation(s):
// \regs[9][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~27_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N9
dffeas \regs[9][19] (
	.clk(CLK),
	.d(\regs[9][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][19] .is_wysiwyg = "true";
defparam \regs[9][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N7
dffeas \regs[11][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][19] .is_wysiwyg = "true";
defparam \regs[11][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N15
dffeas \regs[10][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][19] .is_wysiwyg = "true";
defparam \regs[10][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N16
cycloneive_lcell_comb \Mux44~12 (
// Equation(s):
// \Mux44~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\regs[10][19]~q ))) # (!dcifimemload_17 & (\regs[8][19]~q ))))

	.dataa(\regs[8][19]~q ),
	.datab(\regs[10][19]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux44~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~12 .lut_mask = 16'hFC0A;
defparam \Mux44~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N6
cycloneive_lcell_comb \Mux44~13 (
// Equation(s):
// \Mux44~13_combout  = (dcifimemload_16 & ((\Mux44~12_combout  & ((\regs[11][19]~q ))) # (!\Mux44~12_combout  & (\regs[9][19]~q )))) # (!dcifimemload_16 & (((\Mux44~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][19]~q ),
	.datac(\regs[11][19]~q ),
	.datad(\Mux44~12_combout ),
	.cin(gnd),
	.combout(\Mux44~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~13 .lut_mask = 16'hF588;
defparam \Mux44~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N30
cycloneive_lcell_comb \Mux44~16 (
// Equation(s):
// \Mux44~16_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux44~13_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & (\Mux44~15_combout )))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux44~15_combout ),
	.datad(\Mux44~13_combout ),
	.cin(gnd),
	.combout(\Mux44~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~16 .lut_mask = 16'hBA98;
defparam \Mux44~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N3
dffeas \regs[6][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][19] .is_wysiwyg = "true";
defparam \regs[6][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N24
cycloneive_lcell_comb \regs[7][19]~feeder (
// Equation(s):
// \regs[7][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~27_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[7][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[7][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[7][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N25
dffeas \regs[7][19] (
	.clk(CLK),
	.d(\regs[7][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][19] .is_wysiwyg = "true";
defparam \regs[7][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y45_N25
dffeas \regs[5][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][19] .is_wysiwyg = "true";
defparam \regs[5][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N6
cycloneive_lcell_comb \Mux44~10 (
// Equation(s):
// \Mux44~10_combout  = (dcifimemload_16 & (((\regs[5][19]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][19]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][19]~q ),
	.datab(\regs[5][19]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux44~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~10 .lut_mask = 16'hF0CA;
defparam \Mux44~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N6
cycloneive_lcell_comb \Mux44~11 (
// Equation(s):
// \Mux44~11_combout  = (dcifimemload_17 & ((\Mux44~10_combout  & ((\regs[7][19]~q ))) # (!\Mux44~10_combout  & (\regs[6][19]~q )))) # (!dcifimemload_17 & (((\Mux44~10_combout ))))

	.dataa(\regs[6][19]~q ),
	.datab(\regs[7][19]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux44~10_combout ),
	.cin(gnd),
	.combout(\Mux44~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~11 .lut_mask = 16'hCFA0;
defparam \Mux44~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N5
dffeas \regs[20][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][19] .is_wysiwyg = "true";
defparam \regs[20][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N6
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (dcifimemload_24 & (((\regs[24][19]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[16][19]~q  & ((!dcifimemload_23))))

	.dataa(\regs[16][19]~q ),
	.datab(\regs[24][19]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hF0CA;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N4
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (dcifimemload_23 & ((\Mux12~4_combout  & (\regs[28][19]~q )) # (!\Mux12~4_combout  & ((\regs[20][19]~q ))))) # (!dcifimemload_23 & (((\Mux12~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[28][19]~q ),
	.datac(\regs[20][19]~q ),
	.datad(\Mux12~4_combout ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hDDA0;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N30
cycloneive_lcell_comb \regs[22][19]~feeder (
// Equation(s):
// \regs[22][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~27_combout ),
	.cin(gnd),
	.combout(\regs[22][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[22][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N31
dffeas \regs[22][19] (
	.clk(CLK),
	.d(\regs[22][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][19] .is_wysiwyg = "true";
defparam \regs[22][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N8
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\regs[26][19]~q ))) # (!dcifimemload_24 & (\regs[18][19]~q ))))

	.dataa(dcifimemload_23),
	.datab(\regs[18][19]~q ),
	.datac(\regs[26][19]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hFA44;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N20
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (dcifimemload_23 & ((\Mux12~2_combout  & ((\regs[30][19]~q ))) # (!\Mux12~2_combout  & (\regs[22][19]~q )))) # (!dcifimemload_23 & (((\Mux12~2_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[22][19]~q ),
	.datac(\Mux12~2_combout ),
	.datad(\regs[30][19]~q ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hF858;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N16
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux12~3_combout ))) # (!dcifimemload_22 & (\Mux12~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux12~5_combout ),
	.datad(\Mux12~3_combout ),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hDC98;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N30
cycloneive_lcell_comb \regs[19][19]~feeder (
// Equation(s):
// \regs[19][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~27_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[19][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[19][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N31
dffeas \regs[19][19] (
	.clk(CLK),
	.d(\regs[19][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][19] .is_wysiwyg = "true";
defparam \regs[19][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N22
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (dcifimemload_23 & (((\regs[23][19]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[19][19]~q  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[19][19]~q ),
	.datac(\regs[23][19]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hAAE4;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N12
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// \Mux12~8_combout  = (dcifimemload_24 & ((\Mux12~7_combout  & (\regs[31][19]~q )) # (!\Mux12~7_combout  & ((\regs[27][19]~q ))))) # (!dcifimemload_24 & (((\Mux12~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[31][19]~q ),
	.datac(\Mux12~7_combout ),
	.datad(\regs[27][19]~q ),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hDAD0;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N8
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (dcifimemload_23 & (((\regs[21][19]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[17][19]~q  & ((!dcifimemload_24))))

	.dataa(\regs[17][19]~q ),
	.datab(\regs[21][19]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hF0CA;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N22
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (\Mux12~0_combout  & (((\regs[29][19]~q ) # (!dcifimemload_24)))) # (!\Mux12~0_combout  & (\regs[25][19]~q  & ((dcifimemload_24))))

	.dataa(\regs[25][19]~q ),
	.datab(\regs[29][19]~q ),
	.datac(\Mux12~0_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hCAF0;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N30
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// \Mux12~9_combout  = (dcifimemload_21 & ((\Mux12~6_combout  & (\Mux12~8_combout )) # (!\Mux12~6_combout  & ((\Mux12~1_combout ))))) # (!dcifimemload_21 & (\Mux12~6_combout ))

	.dataa(dcifimemload_21),
	.datab(\Mux12~6_combout ),
	.datac(\Mux12~8_combout ),
	.datad(\Mux12~1_combout ),
	.cin(gnd),
	.combout(\Mux12~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hE6C4;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N14
cycloneive_lcell_comb \Mux12~10 (
// Equation(s):
// \Mux12~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][19]~q ))) # (!dcifimemload_22 & (\regs[8][19]~q ))))

	.dataa(\regs[8][19]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[10][19]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux12~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~10 .lut_mask = 16'hFC22;
defparam \Mux12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N10
cycloneive_lcell_comb \Mux12~11 (
// Equation(s):
// \Mux12~11_combout  = (dcifimemload_21 & ((\Mux12~10_combout  & (\regs[11][19]~q )) # (!\Mux12~10_combout  & ((\regs[9][19]~q ))))) # (!dcifimemload_21 & (((\Mux12~10_combout ))))

	.dataa(\regs[11][19]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[9][19]~q ),
	.datad(\Mux12~10_combout ),
	.cin(gnd),
	.combout(\Mux12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~11 .lut_mask = 16'hBBC0;
defparam \Mux12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N26
cycloneive_lcell_comb \regs[12][19]~feeder (
// Equation(s):
// \regs[12][19]~feeder_combout  = \regs~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~27_combout ),
	.cin(gnd),
	.combout(\regs[12][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[12][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[12][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N27
dffeas \regs[12][19] (
	.clk(CLK),
	.d(\regs[12][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][19] .is_wysiwyg = "true";
defparam \regs[12][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N18
cycloneive_lcell_comb \Mux12~17 (
// Equation(s):
// \Mux12~17_combout  = (dcifimemload_21 & (((\regs[13][19]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][19]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][19]~q ),
	.datac(\regs[13][19]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~17 .lut_mask = 16'hAAE4;
defparam \Mux12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N0
cycloneive_lcell_comb \Mux12~18 (
// Equation(s):
// \Mux12~18_combout  = (dcifimemload_22 & ((\Mux12~17_combout  & (\regs[15][19]~q )) # (!\Mux12~17_combout  & ((\regs[14][19]~q ))))) # (!dcifimemload_22 & (((\Mux12~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][19]~q ),
	.datac(\regs[14][19]~q ),
	.datad(\Mux12~17_combout ),
	.cin(gnd),
	.combout(\Mux12~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~18 .lut_mask = 16'hDDA0;
defparam \Mux12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N9
dffeas \regs[4][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~27_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][19] .is_wysiwyg = "true";
defparam \regs[4][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N24
cycloneive_lcell_comb \Mux12~12 (
// Equation(s):
// \Mux12~12_combout  = (dcifimemload_21 & (((\regs[5][19]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][19]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][19]~q ),
	.datac(\regs[5][19]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~12 .lut_mask = 16'hAAE4;
defparam \Mux12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N2
cycloneive_lcell_comb \Mux12~13 (
// Equation(s):
// \Mux12~13_combout  = (dcifimemload_22 & ((\Mux12~12_combout  & (\regs[7][19]~q )) # (!\Mux12~12_combout  & ((\regs[6][19]~q ))))) # (!dcifimemload_22 & (((\Mux12~12_combout ))))

	.dataa(\regs[7][19]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[6][19]~q ),
	.datad(\Mux12~12_combout ),
	.cin(gnd),
	.combout(\Mux12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~13 .lut_mask = 16'hBBC0;
defparam \Mux12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N16
cycloneive_lcell_comb \Mux12~14 (
// Equation(s):
// \Mux12~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][19]~q ))) # (!dcifimemload_22 & (\regs[1][19]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[1][19]~q ),
	.datac(\regs[3][19]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~14 .lut_mask = 16'hA088;
defparam \Mux12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N12
cycloneive_lcell_comb \Mux12~15 (
// Equation(s):
// \Mux12~15_combout  = (\Mux12~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \regs[2][19]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[2][19]~q ),
	.datad(\Mux12~14_combout ),
	.cin(gnd),
	.combout(\Mux12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~15 .lut_mask = 16'hFF40;
defparam \Mux12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N18
cycloneive_lcell_comb \Mux12~16 (
// Equation(s):
// \Mux12~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux12~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & ((\Mux12~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux12~13_combout ),
	.datad(\Mux12~15_combout ),
	.cin(gnd),
	.combout(\Mux12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~16 .lut_mask = 16'hB9A8;
defparam \Mux12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N28
cycloneive_lcell_comb \Mux12~19 (
// Equation(s):
// \Mux12~19_combout  = (dcifimemload_24 & ((\Mux12~16_combout  & ((\Mux12~18_combout ))) # (!\Mux12~16_combout  & (\Mux12~11_combout )))) # (!dcifimemload_24 & (((\Mux12~16_combout ))))

	.dataa(\Mux12~11_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux12~18_combout ),
	.datad(\Mux12~16_combout ),
	.cin(gnd),
	.combout(\Mux12~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~19 .lut_mask = 16'hF388;
defparam \Mux12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N4
cycloneive_lcell_comb \regs~28 (
// Equation(s):
// \regs~28_combout  = (!\Equal0~1_combout  & \Selector13~1_combout )

	.dataa(\Equal0~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector13),
	.cin(gnd),
	.combout(\regs~28_combout ),
	.cout());
// synopsys translate_off
defparam \regs~28 .lut_mask = 16'h5500;
defparam \regs~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N22
cycloneive_lcell_comb \regs[22][18]~feeder (
// Equation(s):
// \regs[22][18]~feeder_combout  = \regs~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~28_combout ),
	.cin(gnd),
	.combout(\regs[22][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][18]~feeder .lut_mask = 16'hFF00;
defparam \regs[22][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N23
dffeas \regs[22][18] (
	.clk(CLK),
	.d(\regs[22][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][18] .is_wysiwyg = "true";
defparam \regs[22][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N11
dffeas \regs[30][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][18] .is_wysiwyg = "true";
defparam \regs[30][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N1
dffeas \regs[18][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][18] .is_wysiwyg = "true";
defparam \regs[18][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N0
cycloneive_lcell_comb \Mux45~2 (
// Equation(s):
// \Mux45~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[26][18]~q )) # (!dcifimemload_19 & ((\regs[18][18]~q )))))

	.dataa(\regs[26][18]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][18]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux45~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~2 .lut_mask = 16'hEE30;
defparam \Mux45~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N10
cycloneive_lcell_comb \Mux45~3 (
// Equation(s):
// \Mux45~3_combout  = (dcifimemload_18 & ((\Mux45~2_combout  & ((\regs[30][18]~q ))) # (!\Mux45~2_combout  & (\regs[22][18]~q )))) # (!dcifimemload_18 & (((\Mux45~2_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[22][18]~q ),
	.datac(\regs[30][18]~q ),
	.datad(\Mux45~2_combout ),
	.cin(gnd),
	.combout(\Mux45~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~3 .lut_mask = 16'hF588;
defparam \Mux45~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N29
dffeas \regs[20][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][18] .is_wysiwyg = "true";
defparam \regs[20][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N27
dffeas \regs[28][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][18] .is_wysiwyg = "true";
defparam \regs[28][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N26
cycloneive_lcell_comb \Mux45~5 (
// Equation(s):
// \Mux45~5_combout  = (\Mux45~4_combout  & (((\regs[28][18]~q ) # (!dcifimemload_18)))) # (!\Mux45~4_combout  & (\regs[20][18]~q  & ((dcifimemload_18))))

	.dataa(\Mux45~4_combout ),
	.datab(\regs[20][18]~q ),
	.datac(\regs[28][18]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux45~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~5 .lut_mask = 16'hE4AA;
defparam \Mux45~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N4
cycloneive_lcell_comb \Mux45~6 (
// Equation(s):
// \Mux45~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux45~3_combout )) # (!dcifimemload_17 & ((\Mux45~5_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux45~3_combout ),
	.datad(\Mux45~5_combout ),
	.cin(gnd),
	.combout(\Mux45~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~6 .lut_mask = 16'hD9C8;
defparam \Mux45~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N3
dffeas \regs[27][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][18] .is_wysiwyg = "true";
defparam \regs[27][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N29
dffeas \regs[31][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][18] .is_wysiwyg = "true";
defparam \regs[31][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N5
dffeas \regs[23][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][18] .is_wysiwyg = "true";
defparam \regs[23][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N15
dffeas \regs[19][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][18] .is_wysiwyg = "true";
defparam \regs[19][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N14
cycloneive_lcell_comb \Mux45~7 (
// Equation(s):
// \Mux45~7_combout  = (dcifimemload_18 & ((\regs[23][18]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[19][18]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[23][18]~q ),
	.datac(\regs[19][18]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux45~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~7 .lut_mask = 16'hAAD8;
defparam \Mux45~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N28
cycloneive_lcell_comb \Mux45~8 (
// Equation(s):
// \Mux45~8_combout  = (dcifimemload_19 & ((\Mux45~7_combout  & ((\regs[31][18]~q ))) # (!\Mux45~7_combout  & (\regs[27][18]~q )))) # (!dcifimemload_19 & (((\Mux45~7_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[27][18]~q ),
	.datac(\regs[31][18]~q ),
	.datad(\Mux45~7_combout ),
	.cin(gnd),
	.combout(\Mux45~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~8 .lut_mask = 16'hF588;
defparam \Mux45~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N3
dffeas \regs[25][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][18] .is_wysiwyg = "true";
defparam \regs[25][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N13
dffeas \regs[29][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][18] .is_wysiwyg = "true";
defparam \regs[29][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N27
dffeas \regs[21][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][18] .is_wysiwyg = "true";
defparam \regs[21][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N31
dffeas \regs[17][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][18] .is_wysiwyg = "true";
defparam \regs[17][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N30
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[21][18]~q )) # (!dcifimemload_18 & ((\regs[17][18]~q )))))

	.dataa(dcifimemload_19),
	.datab(\regs[21][18]~q ),
	.datac(\regs[17][18]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hEE50;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N12
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (dcifimemload_19 & ((\Mux45~0_combout  & ((\regs[29][18]~q ))) # (!\Mux45~0_combout  & (\regs[25][18]~q )))) # (!dcifimemload_19 & (((\Mux45~0_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[25][18]~q ),
	.datac(\regs[29][18]~q ),
	.datad(\Mux45~0_combout ),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hF588;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N29
dffeas \regs[14][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][18] .is_wysiwyg = "true";
defparam \regs[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N27
dffeas \regs[15][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][18] .is_wysiwyg = "true";
defparam \regs[15][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y43_N7
dffeas \regs[12][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][18] .is_wysiwyg = "true";
defparam \regs[12][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N6
cycloneive_lcell_comb \Mux45~17 (
// Equation(s):
// \Mux45~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][18]~q )) # (!dcifimemload_16 & ((\regs[12][18]~q )))))

	.dataa(\regs[13][18]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][18]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux45~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~17 .lut_mask = 16'hEE30;
defparam \Mux45~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N26
cycloneive_lcell_comb \Mux45~18 (
// Equation(s):
// \Mux45~18_combout  = (dcifimemload_17 & ((\Mux45~17_combout  & ((\regs[15][18]~q ))) # (!\Mux45~17_combout  & (\regs[14][18]~q )))) # (!dcifimemload_17 & (((\Mux45~17_combout ))))

	.dataa(\regs[14][18]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[15][18]~q ),
	.datad(\Mux45~17_combout ),
	.cin(gnd),
	.combout(\Mux45~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~18 .lut_mask = 16'hF388;
defparam \Mux45~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N29
dffeas \regs[9][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][18] .is_wysiwyg = "true";
defparam \regs[9][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N31
dffeas \regs[11][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][18] .is_wysiwyg = "true";
defparam \regs[11][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N21
dffeas \regs[8][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][18] .is_wysiwyg = "true";
defparam \regs[8][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N20
cycloneive_lcell_comb \Mux45~10 (
// Equation(s):
// \Mux45~10_combout  = (dcifimemload_17 & ((\regs[10][18]~q ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((\regs[8][18]~q  & !dcifimemload_16))))

	.dataa(\regs[10][18]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[8][18]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux45~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~10 .lut_mask = 16'hCCB8;
defparam \Mux45~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N30
cycloneive_lcell_comb \Mux45~11 (
// Equation(s):
// \Mux45~11_combout  = (dcifimemload_16 & ((\Mux45~10_combout  & ((\regs[11][18]~q ))) # (!\Mux45~10_combout  & (\regs[9][18]~q )))) # (!dcifimemload_16 & (((\Mux45~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][18]~q ),
	.datac(\regs[11][18]~q ),
	.datad(\Mux45~10_combout ),
	.cin(gnd),
	.combout(\Mux45~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~11 .lut_mask = 16'hF588;
defparam \Mux45~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N25
dffeas \regs[2][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][18] .is_wysiwyg = "true";
defparam \regs[2][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N15
dffeas \regs[1][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][18] .is_wysiwyg = "true";
defparam \regs[1][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N14
cycloneive_lcell_comb \Mux45~14 (
// Equation(s):
// \Mux45~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][18]~q )) # (!dcifimemload_17 & ((\regs[1][18]~q )))))

	.dataa(\regs[3][18]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][18]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux45~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~14 .lut_mask = 16'h88C0;
defparam \Mux45~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N24
cycloneive_lcell_comb \Mux45~15 (
// Equation(s):
// \Mux45~15_combout  = (\Mux45~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][18]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][18]~q ),
	.datad(\Mux45~14_combout ),
	.cin(gnd),
	.combout(\Mux45~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~15 .lut_mask = 16'hFF40;
defparam \Mux45~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N27
dffeas \regs[7][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][18] .is_wysiwyg = "true";
defparam \regs[7][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N12
cycloneive_lcell_comb \regs[5][18]~feeder (
// Equation(s):
// \regs[5][18]~feeder_combout  = \regs~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~28_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[5][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][18]~feeder .lut_mask = 16'hF0F0;
defparam \regs[5][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N13
dffeas \regs[5][18] (
	.clk(CLK),
	.d(\regs[5][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][18] .is_wysiwyg = "true";
defparam \regs[5][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N13
dffeas \regs[4][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][18] .is_wysiwyg = "true";
defparam \regs[4][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N12
cycloneive_lcell_comb \Mux45~12 (
// Equation(s):
// \Mux45~12_combout  = (dcifimemload_16 & ((\regs[5][18]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][18]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[5][18]~q ),
	.datac(\regs[4][18]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux45~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~12 .lut_mask = 16'hAAD8;
defparam \Mux45~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N26
cycloneive_lcell_comb \Mux45~13 (
// Equation(s):
// \Mux45~13_combout  = (dcifimemload_17 & ((\Mux45~12_combout  & ((\regs[7][18]~q ))) # (!\Mux45~12_combout  & (\regs[6][18]~q )))) # (!dcifimemload_17 & (((\Mux45~12_combout ))))

	.dataa(\regs[6][18]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[7][18]~q ),
	.datad(\Mux45~12_combout ),
	.cin(gnd),
	.combout(\Mux45~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~13 .lut_mask = 16'hF388;
defparam \Mux45~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N28
cycloneive_lcell_comb \Mux45~16 (
// Equation(s):
// \Mux45~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux45~13_combout ))) # (!dcifimemload_18 & (\Mux45~15_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux45~15_combout ),
	.datad(\Mux45~13_combout ),
	.cin(gnd),
	.combout(\Mux45~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~16 .lut_mask = 16'hDC98;
defparam \Mux45~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N2
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (dcifimemload_24 & (((\regs[25][18]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[17][18]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[17][18]~q ),
	.datac(\regs[25][18]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hAAE4;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N26
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (dcifimemload_23 & ((\Mux13~0_combout  & (\regs[29][18]~q )) # (!\Mux13~0_combout  & ((\regs[21][18]~q ))))) # (!dcifimemload_23 & (((\Mux13~0_combout ))))

	.dataa(\regs[29][18]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[21][18]~q ),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hBBC0;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N2
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// \Mux13~7_combout  = (dcifimemload_24 & (((\regs[27][18]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[19][18]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[19][18]~q ),
	.datac(\regs[27][18]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hAAE4;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N4
cycloneive_lcell_comb \Mux13~8 (
// Equation(s):
// \Mux13~8_combout  = (dcifimemload_23 & ((\Mux13~7_combout  & (\regs[31][18]~q )) # (!\Mux13~7_combout  & ((\regs[23][18]~q ))))) # (!dcifimemload_23 & (((\Mux13~7_combout ))))

	.dataa(\regs[31][18]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[23][18]~q ),
	.datad(\Mux13~7_combout ),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~8 .lut_mask = 16'hBBC0;
defparam \Mux13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N31
dffeas \regs[24][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][18] .is_wysiwyg = "true";
defparam \regs[24][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N13
dffeas \regs[16][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][18] .is_wysiwyg = "true";
defparam \regs[16][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N28
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[20][18]~q ))) # (!dcifimemload_23 & (\regs[16][18]~q ))))

	.dataa(dcifimemload_24),
	.datab(\regs[16][18]~q ),
	.datac(\regs[20][18]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hFA44;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N30
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// \Mux13~5_combout  = (dcifimemload_24 & ((\Mux13~4_combout  & (\regs[28][18]~q )) # (!\Mux13~4_combout  & ((\regs[24][18]~q ))))) # (!dcifimemload_24 & (((\Mux13~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[28][18]~q ),
	.datac(\regs[24][18]~q ),
	.datad(\Mux13~4_combout ),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hDDA0;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N20
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux13~3_combout )) # (!dcifimemload_22 & ((\Mux13~5_combout )))))

	.dataa(\Mux13~3_combout ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\Mux13~5_combout ),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hE3E0;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N22
cycloneive_lcell_comb \Mux13~9 (
// Equation(s):
// \Mux13~9_combout  = (dcifimemload_21 & ((\Mux13~6_combout  & ((\Mux13~8_combout ))) # (!\Mux13~6_combout  & (\Mux13~1_combout )))) # (!dcifimemload_21 & (((\Mux13~6_combout ))))

	.dataa(\Mux13~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux13~8_combout ),
	.datad(\Mux13~6_combout ),
	.cin(gnd),
	.combout(\Mux13~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~9 .lut_mask = 16'hF388;
defparam \Mux13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N24
cycloneive_lcell_comb \regs[6][18]~feeder (
// Equation(s):
// \regs[6][18]~feeder_combout  = \regs~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~28_combout ),
	.cin(gnd),
	.combout(\regs[6][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][18]~feeder .lut_mask = 16'hFF00;
defparam \regs[6][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N25
dffeas \regs[6][18] (
	.clk(CLK),
	.d(\regs[6][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][18] .is_wysiwyg = "true";
defparam \regs[6][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N28
cycloneive_lcell_comb \Mux13~11 (
// Equation(s):
// \Mux13~11_combout  = (\Mux13~10_combout  & (((\regs[7][18]~q ) # (!dcifimemload_22)))) # (!\Mux13~10_combout  & (\regs[6][18]~q  & (dcifimemload_22)))

	.dataa(\Mux13~10_combout ),
	.datab(\regs[6][18]~q ),
	.datac(dcifimemload_22),
	.datad(\regs[7][18]~q ),
	.cin(gnd),
	.combout(\Mux13~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~11 .lut_mask = 16'hEA4A;
defparam \Mux13~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N28
cycloneive_lcell_comb \Mux13~18 (
// Equation(s):
// \Mux13~18_combout  = (\Mux13~17_combout  & ((\regs[15][18]~q ) # ((!dcifimemload_22)))) # (!\Mux13~17_combout  & (((\regs[14][18]~q  & dcifimemload_22))))

	.dataa(\Mux13~17_combout ),
	.datab(\regs[15][18]~q ),
	.datac(\regs[14][18]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux13~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~18 .lut_mask = 16'hD8AA;
defparam \Mux13~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N4
cycloneive_lcell_comb \Mux13~14 (
// Equation(s):
// \Mux13~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\regs[3][18]~q )) # (!dcifimemload_22 & ((\regs[1][18]~q )))))

	.dataa(\regs[3][18]~q ),
	.datab(\regs[1][18]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux13~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~14 .lut_mask = 16'hA0C0;
defparam \Mux13~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N8
cycloneive_lcell_comb \Mux13~15 (
// Equation(s):
// \Mux13~15_combout  = (\Mux13~14_combout ) # ((\regs[2][18]~q  & (!dcifimemload_21 & dcifimemload_22)))

	.dataa(\regs[2][18]~q ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\Mux13~14_combout ),
	.cin(gnd),
	.combout(\Mux13~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~15 .lut_mask = 16'hFF20;
defparam \Mux13~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N5
dffeas \regs[10][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~28_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][18] .is_wysiwyg = "true";
defparam \regs[10][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \Mux13~12 (
// Equation(s):
// \Mux13~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][18]~q ))) # (!dcifimemload_22 & (\regs[8][18]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][18]~q ),
	.datac(\regs[10][18]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux13~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~12 .lut_mask = 16'hFA44;
defparam \Mux13~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N28
cycloneive_lcell_comb \Mux13~13 (
// Equation(s):
// \Mux13~13_combout  = (dcifimemload_21 & ((\Mux13~12_combout  & (\regs[11][18]~q )) # (!\Mux13~12_combout  & ((\regs[9][18]~q ))))) # (!dcifimemload_21 & (((\Mux13~12_combout ))))

	.dataa(\regs[11][18]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[9][18]~q ),
	.datad(\Mux13~12_combout ),
	.cin(gnd),
	.combout(\Mux13~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~13 .lut_mask = 16'hBBC0;
defparam \Mux13~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N10
cycloneive_lcell_comb \Mux13~16 (
// Equation(s):
// \Mux13~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & ((\Mux13~13_combout ))) # (!dcifimemload_24 & (\Mux13~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux13~15_combout ),
	.datad(\Mux13~13_combout ),
	.cin(gnd),
	.combout(\Mux13~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~16 .lut_mask = 16'hDC98;
defparam \Mux13~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N16
cycloneive_lcell_comb \Mux13~19 (
// Equation(s):
// \Mux13~19_combout  = (dcifimemload_23 & ((\Mux13~16_combout  & ((\Mux13~18_combout ))) # (!\Mux13~16_combout  & (\Mux13~11_combout )))) # (!dcifimemload_23 & (((\Mux13~16_combout ))))

	.dataa(\Mux13~11_combout ),
	.datab(\Mux13~18_combout ),
	.datac(dcifimemload_23),
	.datad(\Mux13~16_combout ),
	.cin(gnd),
	.combout(\Mux13~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~19 .lut_mask = 16'hCFA0;
defparam \Mux13~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N30
cycloneive_lcell_comb \regs~29 (
// Equation(s):
// \regs~29_combout  = (!\Equal0~1_combout  & \Selector14~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Equal0~1_combout ),
	.datad(Selector14),
	.cin(gnd),
	.combout(\regs~29_combout ),
	.cout());
// synopsys translate_off
defparam \regs~29 .lut_mask = 16'h0F00;
defparam \regs~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N31
dffeas \regs[21][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][17] .is_wysiwyg = "true";
defparam \regs[21][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N1
dffeas \regs[29][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][17] .is_wysiwyg = "true";
defparam \regs[29][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N28
cycloneive_lcell_comb \regs[17][17]~feeder (
// Equation(s):
// \regs[17][17]~feeder_combout  = \regs~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~29_combout ),
	.cin(gnd),
	.combout(\regs[17][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][17]~feeder .lut_mask = 16'hFF00;
defparam \regs[17][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N29
dffeas \regs[17][17] (
	.clk(CLK),
	.d(\regs[17][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][17] .is_wysiwyg = "true";
defparam \regs[17][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N6
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (dcifimemload_19 & ((\regs[25][17]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\regs[17][17]~q  & !dcifimemload_18))))

	.dataa(\regs[25][17]~q ),
	.datab(\regs[17][17]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hF0AC;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N0
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (dcifimemload_18 & ((\Mux46~0_combout  & ((\regs[29][17]~q ))) # (!\Mux46~0_combout  & (\regs[21][17]~q )))) # (!dcifimemload_18 & (((\Mux46~0_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[21][17]~q ),
	.datac(\regs[29][17]~q ),
	.datad(\Mux46~0_combout ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hF588;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N27
dffeas \regs[23][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][17] .is_wysiwyg = "true";
defparam \regs[23][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N27
dffeas \regs[31][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][17] .is_wysiwyg = "true";
defparam \regs[31][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N21
dffeas \regs[19][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][17] .is_wysiwyg = "true";
defparam \regs[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N20
cycloneive_lcell_comb \Mux46~7 (
// Equation(s):
// \Mux46~7_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[27][17]~q )) # (!dcifimemload_19 & ((\regs[19][17]~q )))))

	.dataa(\regs[27][17]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[19][17]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux46~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~7 .lut_mask = 16'hEE30;
defparam \Mux46~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N26
cycloneive_lcell_comb \Mux46~8 (
// Equation(s):
// \Mux46~8_combout  = (dcifimemload_18 & ((\Mux46~7_combout  & ((\regs[31][17]~q ))) # (!\Mux46~7_combout  & (\regs[23][17]~q )))) # (!dcifimemload_18 & (((\Mux46~7_combout ))))

	.dataa(\regs[23][17]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[31][17]~q ),
	.datad(\Mux46~7_combout ),
	.cin(gnd),
	.combout(\Mux46~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~8 .lut_mask = 16'hF388;
defparam \Mux46~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N1
dffeas \regs[16][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][17] .is_wysiwyg = "true";
defparam \regs[16][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N0
cycloneive_lcell_comb \Mux46~4 (
// Equation(s):
// \Mux46~4_combout  = (dcifimemload_18 & ((\regs[20][17]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[16][17]~q  & !dcifimemload_19))))

	.dataa(\regs[20][17]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[16][17]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux46~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~4 .lut_mask = 16'hCCB8;
defparam \Mux46~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N7
dffeas \regs[28][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][17] .is_wysiwyg = "true";
defparam \regs[28][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N6
cycloneive_lcell_comb \Mux46~5 (
// Equation(s):
// \Mux46~5_combout  = (\Mux46~4_combout  & (((\regs[28][17]~q ) # (!dcifimemload_19)))) # (!\Mux46~4_combout  & (\regs[24][17]~q  & ((dcifimemload_19))))

	.dataa(\regs[24][17]~q ),
	.datab(\Mux46~4_combout ),
	.datac(\regs[28][17]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux46~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~5 .lut_mask = 16'hE2CC;
defparam \Mux46~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N27
dffeas \regs[30][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][17] .is_wysiwyg = "true";
defparam \regs[30][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N17
dffeas \regs[18][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][17] .is_wysiwyg = "true";
defparam \regs[18][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N16
cycloneive_lcell_comb \Mux46~2 (
// Equation(s):
// \Mux46~2_combout  = (dcifimemload_18 & ((\regs[22][17]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[18][17]~q  & !dcifimemload_19))))

	.dataa(\regs[22][17]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][17]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~2 .lut_mask = 16'hCCB8;
defparam \Mux46~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N26
cycloneive_lcell_comb \Mux46~3 (
// Equation(s):
// \Mux46~3_combout  = (dcifimemload_19 & ((\Mux46~2_combout  & ((\regs[30][17]~q ))) # (!\Mux46~2_combout  & (\regs[26][17]~q )))) # (!dcifimemload_19 & (((\Mux46~2_combout ))))

	.dataa(\regs[26][17]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[30][17]~q ),
	.datad(\Mux46~2_combout ),
	.cin(gnd),
	.combout(\Mux46~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~3 .lut_mask = 16'hF388;
defparam \Mux46~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N16
cycloneive_lcell_comb \Mux46~6 (
// Equation(s):
// \Mux46~6_combout  = (dcifimemload_17 & (((dcifimemload_16) # (\Mux46~3_combout )))) # (!dcifimemload_17 & (\Mux46~5_combout  & (!dcifimemload_16)))

	.dataa(\Mux46~5_combout ),
	.datab(dcifimemload_17),
	.datac(dcifimemload_16),
	.datad(\Mux46~3_combout ),
	.cin(gnd),
	.combout(\Mux46~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~6 .lut_mask = 16'hCEC2;
defparam \Mux46~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N17
dffeas \regs[14][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][17] .is_wysiwyg = "true";
defparam \regs[14][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N9
dffeas \regs[15][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][17] .is_wysiwyg = "true";
defparam \regs[15][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y43_N5
dffeas \regs[12][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][17] .is_wysiwyg = "true";
defparam \regs[12][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N4
cycloneive_lcell_comb \Mux46~17 (
// Equation(s):
// \Mux46~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][17]~q )) # (!dcifimemload_16 & ((\regs[12][17]~q )))))

	.dataa(\regs[13][17]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][17]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux46~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~17 .lut_mask = 16'hEE30;
defparam \Mux46~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N8
cycloneive_lcell_comb \Mux46~18 (
// Equation(s):
// \Mux46~18_combout  = (dcifimemload_17 & ((\Mux46~17_combout  & ((\regs[15][17]~q ))) # (!\Mux46~17_combout  & (\regs[14][17]~q )))) # (!dcifimemload_17 & (((\Mux46~17_combout ))))

	.dataa(\regs[14][17]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[15][17]~q ),
	.datad(\Mux46~17_combout ),
	.cin(gnd),
	.combout(\Mux46~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~18 .lut_mask = 16'hF388;
defparam \Mux46~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N8
cycloneive_lcell_comb \regs[4][17]~feeder (
// Equation(s):
// \regs[4][17]~feeder_combout  = \regs~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~29_combout ),
	.cin(gnd),
	.combout(\regs[4][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[4][17]~feeder .lut_mask = 16'hFF00;
defparam \regs[4][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N9
dffeas \regs[4][17] (
	.clk(CLK),
	.d(\regs[4][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][17] .is_wysiwyg = "true";
defparam \regs[4][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N26
cycloneive_lcell_comb \Mux46~10 (
// Equation(s):
// \Mux46~10_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[5][17]~q )) # (!dcifimemload_16 & ((\regs[4][17]~q )))))

	.dataa(\regs[5][17]~q ),
	.datab(\regs[4][17]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux46~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~10 .lut_mask = 16'hFA0C;
defparam \Mux46~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N9
dffeas \regs[6][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][17] .is_wysiwyg = "true";
defparam \regs[6][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N5
dffeas \regs[7][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][17] .is_wysiwyg = "true";
defparam \regs[7][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N4
cycloneive_lcell_comb \Mux46~11 (
// Equation(s):
// \Mux46~11_combout  = (\Mux46~10_combout  & (((\regs[7][17]~q ) # (!dcifimemload_17)))) # (!\Mux46~10_combout  & (\regs[6][17]~q  & ((dcifimemload_17))))

	.dataa(\Mux46~10_combout ),
	.datab(\regs[6][17]~q ),
	.datac(\regs[7][17]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux46~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~11 .lut_mask = 16'hE4AA;
defparam \Mux46~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N18
cycloneive_lcell_comb \regs[9][17]~feeder (
// Equation(s):
// \regs[9][17]~feeder_combout  = \regs~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~29_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][17]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N19
dffeas \regs[9][17] (
	.clk(CLK),
	.d(\regs[9][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][17] .is_wysiwyg = "true";
defparam \regs[9][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N25
dffeas \regs[10][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][17] .is_wysiwyg = "true";
defparam \regs[10][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N2
cycloneive_lcell_comb \Mux46~12 (
// Equation(s):
// \Mux46~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\regs[10][17]~q ))) # (!dcifimemload_17 & (\regs[8][17]~q ))))

	.dataa(\regs[8][17]~q ),
	.datab(\regs[10][17]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux46~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~12 .lut_mask = 16'hFC0A;
defparam \Mux46~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N14
cycloneive_lcell_comb \Mux46~13 (
// Equation(s):
// \Mux46~13_combout  = (dcifimemload_16 & ((\Mux46~12_combout  & (\regs[11][17]~q )) # (!\Mux46~12_combout  & ((\regs[9][17]~q ))))) # (!dcifimemload_16 & (((\Mux46~12_combout ))))

	.dataa(\regs[11][17]~q ),
	.datab(\regs[9][17]~q ),
	.datac(dcifimemload_16),
	.datad(\Mux46~12_combout ),
	.cin(gnd),
	.combout(\Mux46~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~13 .lut_mask = 16'hAFC0;
defparam \Mux46~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N18
cycloneive_lcell_comb \regs[2][17]~feeder (
// Equation(s):
// \regs[2][17]~feeder_combout  = \regs~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~29_combout ),
	.cin(gnd),
	.combout(\regs[2][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[2][17]~feeder .lut_mask = 16'hFF00;
defparam \regs[2][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N19
dffeas \regs[2][17] (
	.clk(CLK),
	.d(\regs[2][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][17] .is_wysiwyg = "true";
defparam \regs[2][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N23
dffeas \regs[3][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][17] .is_wysiwyg = "true";
defparam \regs[3][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N13
dffeas \regs[1][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][17] .is_wysiwyg = "true";
defparam \regs[1][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N12
cycloneive_lcell_comb \Mux46~14 (
// Equation(s):
// \Mux46~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][17]~q )) # (!dcifimemload_17 & ((\regs[1][17]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[3][17]~q ),
	.datac(\regs[1][17]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux46~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~14 .lut_mask = 16'hD800;
defparam \Mux46~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N2
cycloneive_lcell_comb \Mux46~15 (
// Equation(s):
// \Mux46~15_combout  = (\Mux46~14_combout ) # ((dcifimemload_17 & (\regs[2][17]~q  & !dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\regs[2][17]~q ),
	.datac(dcifimemload_16),
	.datad(\Mux46~14_combout ),
	.cin(gnd),
	.combout(\Mux46~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~15 .lut_mask = 16'hFF08;
defparam \Mux46~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N24
cycloneive_lcell_comb \Mux46~16 (
// Equation(s):
// \Mux46~16_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & (\Mux46~13_combout )) # (!dcifimemload_19 & ((\Mux46~15_combout )))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux46~13_combout ),
	.datad(\Mux46~15_combout ),
	.cin(gnd),
	.combout(\Mux46~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~16 .lut_mask = 16'hD9C8;
defparam \Mux46~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N15
dffeas \regs[27][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][17] .is_wysiwyg = "true";
defparam \regs[27][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N26
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// \Mux14~7_combout  = (dcifimemload_23 & (((\regs[23][17]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[19][17]~q  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[19][17]~q ),
	.datac(\regs[23][17]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'hAAE4;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N14
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (dcifimemload_24 & ((\Mux14~7_combout  & (\regs[31][17]~q )) # (!\Mux14~7_combout  & ((\regs[27][17]~q ))))) # (!dcifimemload_24 & (((\Mux14~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[31][17]~q ),
	.datac(\regs[27][17]~q ),
	.datad(\Mux14~7_combout ),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'hDDA0;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N29
dffeas \regs[20][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][17] .is_wysiwyg = "true";
defparam \regs[20][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N21
dffeas \regs[24][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][17] .is_wysiwyg = "true";
defparam \regs[24][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N20
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[24][17]~q )) # (!dcifimemload_24 & ((\regs[16][17]~q )))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\regs[24][17]~q ),
	.datad(\regs[16][17]~q ),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hD9C8;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N28
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (dcifimemload_23 & ((\Mux14~4_combout  & (\regs[28][17]~q )) # (!\Mux14~4_combout  & ((\regs[20][17]~q ))))) # (!dcifimemload_23 & (((\Mux14~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[28][17]~q ),
	.datac(\regs[20][17]~q ),
	.datad(\Mux14~4_combout ),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hDDA0;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N3
dffeas \regs[22][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][17] .is_wysiwyg = "true";
defparam \regs[22][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N8
cycloneive_lcell_comb \regs[26][17]~feeder (
// Equation(s):
// \regs[26][17]~feeder_combout  = \regs~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~29_combout ),
	.cin(gnd),
	.combout(\regs[26][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][17]~feeder .lut_mask = 16'hFF00;
defparam \regs[26][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N9
dffeas \regs[26][17] (
	.clk(CLK),
	.d(\regs[26][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][17] .is_wysiwyg = "true";
defparam \regs[26][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N10
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\regs[26][17]~q ))) # (!dcifimemload_24 & (\regs[18][17]~q ))))

	.dataa(\regs[18][17]~q ),
	.datab(\regs[26][17]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hFC0A;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N2
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (dcifimemload_23 & ((\Mux14~2_combout  & (\regs[30][17]~q )) # (!\Mux14~2_combout  & ((\regs[22][17]~q ))))) # (!dcifimemload_23 & (((\Mux14~2_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[30][17]~q ),
	.datac(\regs[22][17]~q ),
	.datad(\Mux14~2_combout ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hDDA0;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N26
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// \Mux14~6_combout  = (dcifimemload_22 & (((dcifimemload_21) # (\Mux14~3_combout )))) # (!dcifimemload_22 & (\Mux14~5_combout  & (!dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\Mux14~5_combout ),
	.datac(dcifimemload_21),
	.datad(\Mux14~3_combout ),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hAEA4;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N21
dffeas \regs[25][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][17] .is_wysiwyg = "true";
defparam \regs[25][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N8
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[21][17]~q )) # (!dcifimemload_23 & ((\regs[17][17]~q )))))

	.dataa(\regs[21][17]~q ),
	.datab(\regs[17][17]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hFA0C;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N20
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (dcifimemload_24 & ((\Mux14~0_combout  & (\regs[29][17]~q )) # (!\Mux14~0_combout  & ((\regs[25][17]~q ))))) # (!dcifimemload_24 & (((\Mux14~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[29][17]~q ),
	.datac(\regs[25][17]~q ),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hDDA0;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N12
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// \Mux14~9_combout  = (dcifimemload_21 & ((\Mux14~6_combout  & (\Mux14~8_combout )) # (!\Mux14~6_combout  & ((\Mux14~1_combout ))))) # (!dcifimemload_21 & (((\Mux14~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux14~8_combout ),
	.datac(\Mux14~6_combout ),
	.datad(\Mux14~1_combout ),
	.cin(gnd),
	.combout(\Mux14~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hDAD0;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N24
cycloneive_lcell_comb \Mux14~10 (
// Equation(s):
// \Mux14~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][17]~q ))) # (!dcifimemload_22 & (\regs[8][17]~q ))))

	.dataa(\regs[8][17]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[10][17]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux14~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~10 .lut_mask = 16'hFC22;
defparam \Mux14~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N4
cycloneive_lcell_comb \Mux14~11 (
// Equation(s):
// \Mux14~11_combout  = (dcifimemload_21 & ((\Mux14~10_combout  & (\regs[11][17]~q )) # (!\Mux14~10_combout  & ((\regs[9][17]~q ))))) # (!dcifimemload_21 & (((\Mux14~10_combout ))))

	.dataa(\regs[11][17]~q ),
	.datab(\regs[9][17]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux14~10_combout ),
	.cin(gnd),
	.combout(\Mux14~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~11 .lut_mask = 16'hAFC0;
defparam \Mux14~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N15
dffeas \regs[13][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][17] .is_wysiwyg = "true";
defparam \regs[13][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N14
cycloneive_lcell_comb \Mux14~17 (
// Equation(s):
// \Mux14~17_combout  = (dcifimemload_21 & (((\regs[13][17]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][17]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][17]~q ),
	.datac(\regs[13][17]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux14~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~17 .lut_mask = 16'hAAE4;
defparam \Mux14~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N16
cycloneive_lcell_comb \Mux14~18 (
// Equation(s):
// \Mux14~18_combout  = (dcifimemload_22 & ((\Mux14~17_combout  & ((\regs[15][17]~q ))) # (!\Mux14~17_combout  & (\regs[14][17]~q )))) # (!dcifimemload_22 & (\Mux14~17_combout ))

	.dataa(dcifimemload_22),
	.datab(\Mux14~17_combout ),
	.datac(\regs[14][17]~q ),
	.datad(\regs[15][17]~q ),
	.cin(gnd),
	.combout(\Mux14~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~18 .lut_mask = 16'hEC64;
defparam \Mux14~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N30
cycloneive_lcell_comb \Mux14~14 (
// Equation(s):
// \Mux14~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][17]~q ))) # (!dcifimemload_22 & (\regs[1][17]~q ))))

	.dataa(\regs[1][17]~q ),
	.datab(\regs[3][17]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux14~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~14 .lut_mask = 16'hCA00;
defparam \Mux14~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N28
cycloneive_lcell_comb \Mux14~15 (
// Equation(s):
// \Mux14~15_combout  = (\Mux14~14_combout ) # ((\regs[2][17]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\regs[2][17]~q ),
	.datab(dcifimemload_22),
	.datac(\Mux14~14_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux14~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~15 .lut_mask = 16'hF0F8;
defparam \Mux14~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N1
dffeas \regs[5][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~29_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][17] .is_wysiwyg = "true";
defparam \regs[5][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \Mux14~12 (
// Equation(s):
// \Mux14~12_combout  = (dcifimemload_21 & (((\regs[5][17]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][17]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][17]~q ),
	.datac(\regs[5][17]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux14~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~12 .lut_mask = 16'hAAE4;
defparam \Mux14~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N8
cycloneive_lcell_comb \Mux14~13 (
// Equation(s):
// \Mux14~13_combout  = (dcifimemload_22 & ((\Mux14~12_combout  & (\regs[7][17]~q )) # (!\Mux14~12_combout  & ((\regs[6][17]~q ))))) # (!dcifimemload_22 & (((\Mux14~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[7][17]~q ),
	.datac(\regs[6][17]~q ),
	.datad(\Mux14~12_combout ),
	.cin(gnd),
	.combout(\Mux14~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~13 .lut_mask = 16'hDDA0;
defparam \Mux14~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N18
cycloneive_lcell_comb \Mux14~16 (
// Equation(s):
// \Mux14~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux14~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & (\Mux14~15_combout )))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux14~15_combout ),
	.datad(\Mux14~13_combout ),
	.cin(gnd),
	.combout(\Mux14~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~16 .lut_mask = 16'hBA98;
defparam \Mux14~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N0
cycloneive_lcell_comb \Mux14~19 (
// Equation(s):
// \Mux14~19_combout  = (dcifimemload_24 & ((\Mux14~16_combout  & ((\Mux14~18_combout ))) # (!\Mux14~16_combout  & (\Mux14~11_combout )))) # (!dcifimemload_24 & (((\Mux14~16_combout ))))

	.dataa(\Mux14~11_combout ),
	.datab(\Mux14~18_combout ),
	.datac(dcifimemload_24),
	.datad(\Mux14~16_combout ),
	.cin(gnd),
	.combout(\Mux14~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~19 .lut_mask = 16'hCFA0;
defparam \Mux14~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N22
cycloneive_lcell_comb \regs~30 (
// Equation(s):
// \regs~30_combout  = (!\Equal0~1_combout  & \Selector15~1_combout )

	.dataa(\Equal0~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector15),
	.cin(gnd),
	.combout(\regs~30_combout ),
	.cout());
// synopsys translate_off
defparam \regs~30 .lut_mask = 16'h5500;
defparam \regs~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N23
dffeas \regs[25][16] (
	.clk(CLK),
	.d(\regs~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][16] .is_wysiwyg = "true";
defparam \regs[25][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N5
dffeas \regs[29][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][16] .is_wysiwyg = "true";
defparam \regs[29][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N18
cycloneive_lcell_comb \regs[21][16]~feeder (
// Equation(s):
// \regs[21][16]~feeder_combout  = \regs~30_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~30_combout ),
	.cin(gnd),
	.combout(\regs[21][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][16]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N19
dffeas \regs[21][16] (
	.clk(CLK),
	.d(\regs[21][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][16] .is_wysiwyg = "true";
defparam \regs[21][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N19
dffeas \regs[17][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][16] .is_wysiwyg = "true";
defparam \regs[17][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N18
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (dcifimemload_18 & ((\regs[21][16]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[17][16]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[21][16]~q ),
	.datac(\regs[17][16]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hAAD8;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N4
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (dcifimemload_19 & ((\Mux47~0_combout  & ((\regs[29][16]~q ))) # (!\Mux47~0_combout  & (\regs[25][16]~q )))) # (!dcifimemload_19 & (((\Mux47~0_combout ))))

	.dataa(\regs[25][16]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[29][16]~q ),
	.datad(\Mux47~0_combout ),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hF388;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N14
cycloneive_lcell_comb \regs[22][16]~feeder (
// Equation(s):
// \regs[22][16]~feeder_combout  = \regs~30_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~30_combout ),
	.cin(gnd),
	.combout(\regs[22][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[22][16]~feeder .lut_mask = 16'hFF00;
defparam \regs[22][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N15
dffeas \regs[22][16] (
	.clk(CLK),
	.d(\regs[22][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][16] .is_wysiwyg = "true";
defparam \regs[22][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N7
dffeas \regs[30][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][16] .is_wysiwyg = "true";
defparam \regs[30][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N29
dffeas \regs[18][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][16] .is_wysiwyg = "true";
defparam \regs[18][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N28
cycloneive_lcell_comb \Mux47~2 (
// Equation(s):
// \Mux47~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[26][16]~q )) # (!dcifimemload_19 & ((\regs[18][16]~q )))))

	.dataa(\regs[26][16]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][16]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux47~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~2 .lut_mask = 16'hEE30;
defparam \Mux47~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N6
cycloneive_lcell_comb \Mux47~3 (
// Equation(s):
// \Mux47~3_combout  = (dcifimemload_18 & ((\Mux47~2_combout  & ((\regs[30][16]~q ))) # (!\Mux47~2_combout  & (\regs[22][16]~q )))) # (!dcifimemload_18 & (((\Mux47~2_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[22][16]~q ),
	.datac(\regs[30][16]~q ),
	.datad(\Mux47~2_combout ),
	.cin(gnd),
	.combout(\Mux47~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~3 .lut_mask = 16'hF588;
defparam \Mux47~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N5
dffeas \regs[20][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][16] .is_wysiwyg = "true";
defparam \regs[20][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N19
dffeas \regs[28][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][16] .is_wysiwyg = "true";
defparam \regs[28][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N28
cycloneive_lcell_comb \regs[24][16]~feeder (
// Equation(s):
// \regs[24][16]~feeder_combout  = \regs~30_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~30_combout ),
	.cin(gnd),
	.combout(\regs[24][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][16]~feeder .lut_mask = 16'hFF00;
defparam \regs[24][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N29
dffeas \regs[24][16] (
	.clk(CLK),
	.d(\regs[24][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][16] .is_wysiwyg = "true";
defparam \regs[24][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N25
dffeas \regs[16][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][16] .is_wysiwyg = "true";
defparam \regs[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N24
cycloneive_lcell_comb \Mux47~4 (
// Equation(s):
// \Mux47~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[24][16]~q )) # (!dcifimemload_19 & ((\regs[16][16]~q )))))

	.dataa(dcifimemload_18),
	.datab(\regs[24][16]~q ),
	.datac(\regs[16][16]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux47~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~4 .lut_mask = 16'hEE50;
defparam \Mux47~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N18
cycloneive_lcell_comb \Mux47~5 (
// Equation(s):
// \Mux47~5_combout  = (dcifimemload_18 & ((\Mux47~4_combout  & ((\regs[28][16]~q ))) # (!\Mux47~4_combout  & (\regs[20][16]~q )))) # (!dcifimemload_18 & (((\Mux47~4_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[20][16]~q ),
	.datac(\regs[28][16]~q ),
	.datad(\Mux47~4_combout ),
	.cin(gnd),
	.combout(\Mux47~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~5 .lut_mask = 16'hF588;
defparam \Mux47~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N20
cycloneive_lcell_comb \Mux47~6 (
// Equation(s):
// \Mux47~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux47~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & ((\Mux47~5_combout ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux47~3_combout ),
	.datad(\Mux47~5_combout ),
	.cin(gnd),
	.combout(\Mux47~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~6 .lut_mask = 16'hB9A8;
defparam \Mux47~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N26
cycloneive_lcell_comb \regs[27][16]~feeder (
// Equation(s):
// \regs[27][16]~feeder_combout  = \regs~30_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~30_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][16]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N27
dffeas \regs[27][16] (
	.clk(CLK),
	.d(\regs[27][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][16] .is_wysiwyg = "true";
defparam \regs[27][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N13
dffeas \regs[31][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][16] .is_wysiwyg = "true";
defparam \regs[31][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N9
dffeas \regs[23][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][16] .is_wysiwyg = "true";
defparam \regs[23][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N23
dffeas \regs[19][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][16] .is_wysiwyg = "true";
defparam \regs[19][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N22
cycloneive_lcell_comb \Mux47~7 (
// Equation(s):
// \Mux47~7_combout  = (dcifimemload_18 & ((\regs[23][16]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[19][16]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[23][16]~q ),
	.datac(\regs[19][16]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux47~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~7 .lut_mask = 16'hAAD8;
defparam \Mux47~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N12
cycloneive_lcell_comb \Mux47~8 (
// Equation(s):
// \Mux47~8_combout  = (dcifimemload_19 & ((\Mux47~7_combout  & ((\regs[31][16]~q ))) # (!\Mux47~7_combout  & (\regs[27][16]~q )))) # (!dcifimemload_19 & (((\Mux47~7_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[27][16]~q ),
	.datac(\regs[31][16]~q ),
	.datad(\Mux47~7_combout ),
	.cin(gnd),
	.combout(\Mux47~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~8 .lut_mask = 16'hF588;
defparam \Mux47~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N25
dffeas \regs[14][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][16] .is_wysiwyg = "true";
defparam \regs[14][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N22
cycloneive_lcell_comb \regs[15][16]~feeder (
// Equation(s):
// \regs[15][16]~feeder_combout  = \regs~30_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~30_combout ),
	.cin(gnd),
	.combout(\regs[15][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][16]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N23
dffeas \regs[15][16] (
	.clk(CLK),
	.d(\regs[15][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][16] .is_wysiwyg = "true";
defparam \regs[15][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y43_N3
dffeas \regs[12][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][16] .is_wysiwyg = "true";
defparam \regs[12][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N2
cycloneive_lcell_comb \Mux47~17 (
// Equation(s):
// \Mux47~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][16]~q )) # (!dcifimemload_16 & ((\regs[12][16]~q )))))

	.dataa(\regs[13][16]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][16]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux47~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~17 .lut_mask = 16'hEE30;
defparam \Mux47~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N20
cycloneive_lcell_comb \Mux47~18 (
// Equation(s):
// \Mux47~18_combout  = (dcifimemload_17 & ((\Mux47~17_combout  & ((\regs[15][16]~q ))) # (!\Mux47~17_combout  & (\regs[14][16]~q )))) # (!dcifimemload_17 & (((\Mux47~17_combout ))))

	.dataa(\regs[14][16]~q ),
	.datab(\regs[15][16]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux47~17_combout ),
	.cin(gnd),
	.combout(\Mux47~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~18 .lut_mask = 16'hCFA0;
defparam \Mux47~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N14
cycloneive_lcell_comb \regs[9][16]~feeder (
// Equation(s):
// \regs[9][16]~feeder_combout  = \regs~30_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~30_combout ),
	.cin(gnd),
	.combout(\regs[9][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][16]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N15
dffeas \regs[9][16] (
	.clk(CLK),
	.d(\regs[9][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][16] .is_wysiwyg = "true";
defparam \regs[9][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N11
dffeas \regs[11][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][16] .is_wysiwyg = "true";
defparam \regs[11][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N27
dffeas \regs[10][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][16] .is_wysiwyg = "true";
defparam \regs[10][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N25
dffeas \regs[8][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][16] .is_wysiwyg = "true";
defparam \regs[8][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N24
cycloneive_lcell_comb \Mux47~10 (
// Equation(s):
// \Mux47~10_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][16]~q )) # (!dcifimemload_17 & ((\regs[8][16]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][16]~q ),
	.datac(\regs[8][16]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux47~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~10 .lut_mask = 16'hEE50;
defparam \Mux47~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N10
cycloneive_lcell_comb \Mux47~11 (
// Equation(s):
// \Mux47~11_combout  = (dcifimemload_16 & ((\Mux47~10_combout  & ((\regs[11][16]~q ))) # (!\Mux47~10_combout  & (\regs[9][16]~q )))) # (!dcifimemload_16 & (((\Mux47~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][16]~q ),
	.datac(\regs[11][16]~q ),
	.datad(\Mux47~10_combout ),
	.cin(gnd),
	.combout(\Mux47~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~11 .lut_mask = 16'hF588;
defparam \Mux47~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N1
dffeas \regs[2][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][16] .is_wysiwyg = "true";
defparam \regs[2][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N31
dffeas \regs[1][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][16] .is_wysiwyg = "true";
defparam \regs[1][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N30
cycloneive_lcell_comb \Mux47~14 (
// Equation(s):
// \Mux47~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][16]~q )) # (!dcifimemload_17 & ((\regs[1][16]~q )))))

	.dataa(\regs[3][16]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[1][16]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux47~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~14 .lut_mask = 16'hB800;
defparam \Mux47~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N26
cycloneive_lcell_comb \Mux47~15 (
// Equation(s):
// \Mux47~15_combout  = (\Mux47~14_combout ) # ((!dcifimemload_16 & (\regs[2][16]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\regs[2][16]~q ),
	.datac(\Mux47~14_combout ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux47~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~15 .lut_mask = 16'hF4F0;
defparam \Mux47~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N3
dffeas \regs[6][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][16] .is_wysiwyg = "true";
defparam \regs[6][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N29
dffeas \regs[7][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][16] .is_wysiwyg = "true";
defparam \regs[7][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N25
dffeas \regs[5][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][16] .is_wysiwyg = "true";
defparam \regs[5][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N19
dffeas \regs[4][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][16] .is_wysiwyg = "true";
defparam \regs[4][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N18
cycloneive_lcell_comb \Mux47~12 (
// Equation(s):
// \Mux47~12_combout  = (dcifimemload_16 & ((\regs[5][16]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][16]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[5][16]~q ),
	.datac(\regs[4][16]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux47~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~12 .lut_mask = 16'hAAD8;
defparam \Mux47~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N28
cycloneive_lcell_comb \Mux47~13 (
// Equation(s):
// \Mux47~13_combout  = (dcifimemload_17 & ((\Mux47~12_combout  & ((\regs[7][16]~q ))) # (!\Mux47~12_combout  & (\regs[6][16]~q )))) # (!dcifimemload_17 & (((\Mux47~12_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][16]~q ),
	.datac(\regs[7][16]~q ),
	.datad(\Mux47~12_combout ),
	.cin(gnd),
	.combout(\Mux47~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~13 .lut_mask = 16'hF588;
defparam \Mux47~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N28
cycloneive_lcell_comb \Mux47~16 (
// Equation(s):
// \Mux47~16_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux47~13_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & (\Mux47~15_combout )))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux47~15_combout ),
	.datad(\Mux47~13_combout ),
	.cin(gnd),
	.combout(\Mux47~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~16 .lut_mask = 16'hBA98;
defparam \Mux47~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N3
dffeas \regs[13][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][16] .is_wysiwyg = "true";
defparam \regs[13][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N2
cycloneive_lcell_comb \Mux15~17 (
// Equation(s):
// \Mux15~17_combout  = (dcifimemload_21 & (((\regs[13][16]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][16]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][16]~q ),
	.datac(\regs[13][16]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux15~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~17 .lut_mask = 16'hAAE4;
defparam \Mux15~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N24
cycloneive_lcell_comb \Mux15~18 (
// Equation(s):
// \Mux15~18_combout  = (dcifimemload_22 & ((\Mux15~17_combout  & (\regs[15][16]~q )) # (!\Mux15~17_combout  & ((\regs[14][16]~q ))))) # (!dcifimemload_22 & (((\Mux15~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][16]~q ),
	.datac(\regs[14][16]~q ),
	.datad(\Mux15~17_combout ),
	.cin(gnd),
	.combout(\Mux15~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~18 .lut_mask = 16'hDDA0;
defparam \Mux15~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N24
cycloneive_lcell_comb \Mux15~10 (
// Equation(s):
// \Mux15~10_combout  = (dcifimemload_21 & (((\regs[5][16]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][16]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][16]~q ),
	.datac(\regs[5][16]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~10 .lut_mask = 16'hAAE4;
defparam \Mux15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N2
cycloneive_lcell_comb \Mux15~11 (
// Equation(s):
// \Mux15~11_combout  = (dcifimemload_22 & ((\Mux15~10_combout  & (\regs[7][16]~q )) # (!\Mux15~10_combout  & ((\regs[6][16]~q ))))) # (!dcifimemload_22 & (((\Mux15~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[7][16]~q ),
	.datac(\regs[6][16]~q ),
	.datad(\Mux15~10_combout ),
	.cin(gnd),
	.combout(\Mux15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~11 .lut_mask = 16'hDDA0;
defparam \Mux15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N13
dffeas \regs[3][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][16] .is_wysiwyg = "true";
defparam \regs[3][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N12
cycloneive_lcell_comb \Mux15~14 (
// Equation(s):
// \Mux15~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][16]~q ))) # (!dcifimemload_22 & (\regs[1][16]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[1][16]~q ),
	.datac(\regs[3][16]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux15~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~14 .lut_mask = 16'hA088;
defparam \Mux15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N28
cycloneive_lcell_comb \Mux15~15 (
// Equation(s):
// \Mux15~15_combout  = (\Mux15~14_combout ) # ((dcifimemload_22 & (\regs[2][16]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\regs[2][16]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux15~14_combout ),
	.cin(gnd),
	.combout(\Mux15~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~15 .lut_mask = 16'hFF08;
defparam \Mux15~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \Mux15~12 (
// Equation(s):
// \Mux15~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][16]~q ))) # (!dcifimemload_22 & (\regs[8][16]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][16]~q ),
	.datac(\regs[10][16]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~12 .lut_mask = 16'hFA44;
defparam \Mux15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N4
cycloneive_lcell_comb \Mux15~13 (
// Equation(s):
// \Mux15~13_combout  = (dcifimemload_21 & ((\Mux15~12_combout  & (\regs[11][16]~q )) # (!\Mux15~12_combout  & ((\regs[9][16]~q ))))) # (!dcifimemload_21 & (((\Mux15~12_combout ))))

	.dataa(\regs[11][16]~q ),
	.datab(\regs[9][16]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux15~12_combout ),
	.cin(gnd),
	.combout(\Mux15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~13 .lut_mask = 16'hAFC0;
defparam \Mux15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N6
cycloneive_lcell_comb \Mux15~16 (
// Equation(s):
// \Mux15~16_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\Mux15~13_combout ))) # (!dcifimemload_24 & (\Mux15~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux15~15_combout ),
	.datac(dcifimemload_24),
	.datad(\Mux15~13_combout ),
	.cin(gnd),
	.combout(\Mux15~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~16 .lut_mask = 16'hF4A4;
defparam \Mux15~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N8
cycloneive_lcell_comb \Mux15~19 (
// Equation(s):
// \Mux15~19_combout  = (dcifimemload_23 & ((\Mux15~16_combout  & (\Mux15~18_combout )) # (!\Mux15~16_combout  & ((\Mux15~11_combout ))))) # (!dcifimemload_23 & (((\Mux15~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux15~18_combout ),
	.datac(\Mux15~11_combout ),
	.datad(\Mux15~16_combout ),
	.cin(gnd),
	.combout(\Mux15~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~19 .lut_mask = 16'hDDA0;
defparam \Mux15~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N12
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// \Mux15~7_combout  = (dcifimemload_24 & ((\regs[27][16]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[19][16]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][16]~q ),
	.datac(\regs[19][16]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'hAAD8;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N8
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// \Mux15~8_combout  = (dcifimemload_23 & ((\Mux15~7_combout  & (\regs[31][16]~q )) # (!\Mux15~7_combout  & ((\regs[23][16]~q ))))) # (!dcifimemload_23 & (((\Mux15~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[31][16]~q ),
	.datac(\regs[23][16]~q ),
	.datad(\Mux15~7_combout ),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hDDA0;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N24
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (dcifimemload_24 & (((dcifimemload_23) # (\regs[25][16]~q )))) # (!dcifimemload_24 & (\regs[17][16]~q  & (!dcifimemload_23)))

	.dataa(dcifimemload_24),
	.datab(\regs[17][16]~q ),
	.datac(dcifimemload_23),
	.datad(\regs[25][16]~q ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hAEA4;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N10
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (dcifimemload_23 & ((\Mux15~0_combout  & (\regs[29][16]~q )) # (!\Mux15~0_combout  & ((\regs[21][16]~q ))))) # (!dcifimemload_23 & (((\Mux15~0_combout ))))

	.dataa(\regs[29][16]~q ),
	.datab(\regs[21][16]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hAFC0;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N4
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[20][16]~q ))) # (!dcifimemload_23 & (\regs[16][16]~q ))))

	.dataa(dcifimemload_24),
	.datab(\regs[16][16]~q ),
	.datac(\regs[20][16]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hFA44;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N26
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (\Mux15~4_combout  & ((\regs[28][16]~q ) # ((!dcifimemload_24)))) # (!\Mux15~4_combout  & (((\regs[24][16]~q  & dcifimemload_24))))

	.dataa(\regs[28][16]~q ),
	.datab(\regs[24][16]~q ),
	.datac(\Mux15~4_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hACF0;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N21
dffeas \regs[26][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~30_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][16] .is_wysiwyg = "true";
defparam \regs[26][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N0
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (dcifimemload_23 & (((\regs[22][16]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[18][16]~q  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[18][16]~q ),
	.datac(\regs[22][16]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hAAE4;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N20
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (dcifimemload_24 & ((\Mux15~2_combout  & (\regs[30][16]~q )) # (!\Mux15~2_combout  & ((\regs[26][16]~q ))))) # (!dcifimemload_24 & (((\Mux15~2_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[30][16]~q ),
	.datac(\regs[26][16]~q ),
	.datad(\Mux15~2_combout ),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hDDA0;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N20
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// \Mux15~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux15~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux15~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux15~5_combout ),
	.datad(\Mux15~3_combout ),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hBA98;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N2
cycloneive_lcell_comb \Mux15~9 (
// Equation(s):
// \Mux15~9_combout  = (dcifimemload_21 & ((\Mux15~6_combout  & (\Mux15~8_combout )) # (!\Mux15~6_combout  & ((\Mux15~1_combout ))))) # (!dcifimemload_21 & (((\Mux15~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux15~8_combout ),
	.datac(\Mux15~1_combout ),
	.datad(\Mux15~6_combout ),
	.cin(gnd),
	.combout(\Mux15~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~9 .lut_mask = 16'hDDA0;
defparam \Mux15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N30
cycloneive_lcell_comb \regs~31 (
// Equation(s):
// \regs~31_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_15)) # (!cuifRegSel_0 & ((Mux163)))))

	.dataa(cuifRegSel_0),
	.datab(ramiframload_15),
	.datac(cuifRegSel_11),
	.datad(Mux161),
	.cin(gnd),
	.combout(\regs~31_combout ),
	.cout());
// synopsys translate_off
defparam \regs~31 .lut_mask = 16'h0D08;
defparam \regs~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N8
cycloneive_lcell_comb \regs~32 (
// Equation(s):
// \regs~32_combout  = (!\Equal0~1_combout  & ((\regs~31_combout ) # ((\regs~64_combout  & \Add1~26_combout ))))

	.dataa(\regs~64_combout ),
	.datab(Add113),
	.datac(\regs~31_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\regs~32_combout ),
	.cout());
// synopsys translate_off
defparam \regs~32 .lut_mask = 16'h00F8;
defparam \regs~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N17
dffeas \regs[26][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][15] .is_wysiwyg = "true";
defparam \regs[26][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N3
dffeas \regs[30][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][15] .is_wysiwyg = "true";
defparam \regs[30][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N17
dffeas \regs[22][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][15] .is_wysiwyg = "true";
defparam \regs[22][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N13
dffeas \regs[18][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][15] .is_wysiwyg = "true";
defparam \regs[18][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N12
cycloneive_lcell_comb \Mux48~2 (
// Equation(s):
// \Mux48~2_combout  = (dcifimemload_18 & ((\regs[22][15]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[18][15]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[22][15]~q ),
	.datac(\regs[18][15]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~2 .lut_mask = 16'hAAD8;
defparam \Mux48~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N2
cycloneive_lcell_comb \Mux48~3 (
// Equation(s):
// \Mux48~3_combout  = (dcifimemload_19 & ((\Mux48~2_combout  & ((\regs[30][15]~q ))) # (!\Mux48~2_combout  & (\regs[26][15]~q )))) # (!dcifimemload_19 & (((\Mux48~2_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[26][15]~q ),
	.datac(\regs[30][15]~q ),
	.datad(\Mux48~2_combout ),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~3 .lut_mask = 16'hF588;
defparam \Mux48~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N3
dffeas \regs[20][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][15] .is_wysiwyg = "true";
defparam \regs[20][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N22
cycloneive_lcell_comb \regs[16][15]~feeder (
// Equation(s):
// \regs[16][15]~feeder_combout  = \regs~32_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~32_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[16][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[16][15]~feeder .lut_mask = 16'hF0F0;
defparam \regs[16][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N23
dffeas \regs[16][15] (
	.clk(CLK),
	.d(\regs[16][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][15] .is_wysiwyg = "true";
defparam \regs[16][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N8
cycloneive_lcell_comb \Mux48~4 (
// Equation(s):
// \Mux48~4_combout  = (dcifimemload_18 & ((\regs[20][15]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[16][15]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[20][15]~q ),
	.datac(\regs[16][15]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~4 .lut_mask = 16'hAAD8;
defparam \Mux48~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N15
dffeas \regs[28][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][15] .is_wysiwyg = "true";
defparam \regs[28][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N14
cycloneive_lcell_comb \Mux48~5 (
// Equation(s):
// \Mux48~5_combout  = (\Mux48~4_combout  & (((\regs[28][15]~q ) # (!dcifimemload_19)))) # (!\Mux48~4_combout  & (\regs[24][15]~q  & ((dcifimemload_19))))

	.dataa(\regs[24][15]~q ),
	.datab(\Mux48~4_combout ),
	.datac(\regs[28][15]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~5 .lut_mask = 16'hE2CC;
defparam \Mux48~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N10
cycloneive_lcell_comb \Mux48~6 (
// Equation(s):
// \Mux48~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux48~3_combout )) # (!dcifimemload_17 & ((\Mux48~5_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux48~3_combout ),
	.datad(\Mux48~5_combout ),
	.cin(gnd),
	.combout(\Mux48~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~6 .lut_mask = 16'hD9C8;
defparam \Mux48~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N19
dffeas \regs[21][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][15] .is_wysiwyg = "true";
defparam \regs[21][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N11
dffeas \regs[29][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][15] .is_wysiwyg = "true";
defparam \regs[29][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N28
cycloneive_lcell_comb \regs[25][15]~feeder (
// Equation(s):
// \regs[25][15]~feeder_combout  = \regs~32_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~32_combout ),
	.cin(gnd),
	.combout(\regs[25][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[25][15]~feeder .lut_mask = 16'hFF00;
defparam \regs[25][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N29
dffeas \regs[25][15] (
	.clk(CLK),
	.d(\regs[25][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][15] .is_wysiwyg = "true";
defparam \regs[25][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N10
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (dcifimemload_19 & (((\regs[25][15]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\regs[17][15]~q  & ((!dcifimemload_18))))

	.dataa(\regs[17][15]~q ),
	.datab(\regs[25][15]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hF0CA;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N10
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (dcifimemload_18 & ((\Mux48~0_combout  & ((\regs[29][15]~q ))) # (!\Mux48~0_combout  & (\regs[21][15]~q )))) # (!dcifimemload_18 & (((\Mux48~0_combout ))))

	.dataa(\regs[21][15]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[29][15]~q ),
	.datad(\Mux48~0_combout ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hF388;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N31
dffeas \regs[23][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][15] .is_wysiwyg = "true";
defparam \regs[23][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N19
dffeas \regs[31][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][15] .is_wysiwyg = "true";
defparam \regs[31][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N28
cycloneive_lcell_comb \regs[27][15]~feeder (
// Equation(s):
// \regs[27][15]~feeder_combout  = \regs~32_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~32_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][15]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N29
dffeas \regs[27][15] (
	.clk(CLK),
	.d(\regs[27][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][15] .is_wysiwyg = "true";
defparam \regs[27][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N31
dffeas \regs[19][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][15] .is_wysiwyg = "true";
defparam \regs[19][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N30
cycloneive_lcell_comb \Mux48~7 (
// Equation(s):
// \Mux48~7_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[27][15]~q )) # (!dcifimemload_19 & ((\regs[19][15]~q )))))

	.dataa(dcifimemload_18),
	.datab(\regs[27][15]~q ),
	.datac(\regs[19][15]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux48~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~7 .lut_mask = 16'hEE50;
defparam \Mux48~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N18
cycloneive_lcell_comb \Mux48~8 (
// Equation(s):
// \Mux48~8_combout  = (dcifimemload_18 & ((\Mux48~7_combout  & ((\regs[31][15]~q ))) # (!\Mux48~7_combout  & (\regs[23][15]~q )))) # (!dcifimemload_18 & (((\Mux48~7_combout ))))

	.dataa(\regs[23][15]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[31][15]~q ),
	.datad(\Mux48~7_combout ),
	.cin(gnd),
	.combout(\Mux48~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~8 .lut_mask = 16'hF388;
defparam \Mux48~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N7
dffeas \regs[6][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][15] .is_wysiwyg = "true";
defparam \regs[6][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N25
dffeas \regs[7][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][15] .is_wysiwyg = "true";
defparam \regs[7][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N3
dffeas \regs[4][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][15] .is_wysiwyg = "true";
defparam \regs[4][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N21
dffeas \regs[5][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][15] .is_wysiwyg = "true";
defparam \regs[5][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N2
cycloneive_lcell_comb \Mux48~10 (
// Equation(s):
// \Mux48~10_combout  = (dcifimemload_16 & ((dcifimemload_17) # ((\regs[5][15]~q )))) # (!dcifimemload_16 & (!dcifimemload_17 & (\regs[4][15]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[4][15]~q ),
	.datad(\regs[5][15]~q ),
	.cin(gnd),
	.combout(\Mux48~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~10 .lut_mask = 16'hBA98;
defparam \Mux48~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N24
cycloneive_lcell_comb \Mux48~11 (
// Equation(s):
// \Mux48~11_combout  = (dcifimemload_17 & ((\Mux48~10_combout  & ((\regs[7][15]~q ))) # (!\Mux48~10_combout  & (\regs[6][15]~q )))) # (!dcifimemload_17 & (((\Mux48~10_combout ))))

	.dataa(\regs[6][15]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[7][15]~q ),
	.datad(\Mux48~10_combout ),
	.cin(gnd),
	.combout(\Mux48~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~11 .lut_mask = 16'hF388;
defparam \Mux48~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N12
cycloneive_lcell_comb \regs[15][15]~feeder (
// Equation(s):
// \regs[15][15]~feeder_combout  = \regs~32_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~32_combout ),
	.cin(gnd),
	.combout(\regs[15][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][15]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N13
dffeas \regs[15][15] (
	.clk(CLK),
	.d(\regs[15][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][15] .is_wysiwyg = "true";
defparam \regs[15][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N21
dffeas \regs[14][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][15] .is_wysiwyg = "true";
defparam \regs[14][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y43_N31
dffeas \regs[12][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][15] .is_wysiwyg = "true";
defparam \regs[12][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N30
cycloneive_lcell_comb \Mux48~17 (
// Equation(s):
// \Mux48~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][15]~q )) # (!dcifimemload_16 & ((\regs[12][15]~q )))))

	.dataa(\regs[13][15]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][15]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux48~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~17 .lut_mask = 16'hEE30;
defparam \Mux48~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N22
cycloneive_lcell_comb \Mux48~18 (
// Equation(s):
// \Mux48~18_combout  = (\Mux48~17_combout  & ((\regs[15][15]~q ) # ((!dcifimemload_17)))) # (!\Mux48~17_combout  & (((\regs[14][15]~q  & dcifimemload_17))))

	.dataa(\regs[15][15]~q ),
	.datab(\regs[14][15]~q ),
	.datac(\Mux48~17_combout ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux48~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~18 .lut_mask = 16'hACF0;
defparam \Mux48~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N3
dffeas \regs[2][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][15] .is_wysiwyg = "true";
defparam \regs[2][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N11
dffeas \regs[1][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][15] .is_wysiwyg = "true";
defparam \regs[1][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N10
cycloneive_lcell_comb \Mux48~14 (
// Equation(s):
// \Mux48~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][15]~q )) # (!dcifimemload_17 & ((\regs[1][15]~q )))))

	.dataa(\regs[3][15]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[1][15]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux48~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~14 .lut_mask = 16'hB800;
defparam \Mux48~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N2
cycloneive_lcell_comb \Mux48~15 (
// Equation(s):
// \Mux48~15_combout  = (\Mux48~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][15]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][15]~q ),
	.datad(\Mux48~14_combout ),
	.cin(gnd),
	.combout(\Mux48~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~15 .lut_mask = 16'hFF40;
defparam \Mux48~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N14
cycloneive_lcell_comb \regs[9][15]~feeder (
// Equation(s):
// \regs[9][15]~feeder_combout  = \regs~32_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~32_combout ),
	.cin(gnd),
	.combout(\regs[9][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][15]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N15
dffeas \regs[9][15] (
	.clk(CLK),
	.d(\regs[9][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][15] .is_wysiwyg = "true";
defparam \regs[9][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N23
dffeas \regs[11][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][15] .is_wysiwyg = "true";
defparam \regs[11][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N29
dffeas \regs[8][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][15] .is_wysiwyg = "true";
defparam \regs[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N28
cycloneive_lcell_comb \Mux48~12 (
// Equation(s):
// \Mux48~12_combout  = (dcifimemload_17 & ((\regs[10][15]~q ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((\regs[8][15]~q  & !dcifimemload_16))))

	.dataa(\regs[10][15]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[8][15]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux48~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~12 .lut_mask = 16'hCCB8;
defparam \Mux48~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N22
cycloneive_lcell_comb \Mux48~13 (
// Equation(s):
// \Mux48~13_combout  = (dcifimemload_16 & ((\Mux48~12_combout  & ((\regs[11][15]~q ))) # (!\Mux48~12_combout  & (\regs[9][15]~q )))) # (!dcifimemload_16 & (((\Mux48~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][15]~q ),
	.datac(\regs[11][15]~q ),
	.datad(\Mux48~12_combout ),
	.cin(gnd),
	.combout(\Mux48~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~13 .lut_mask = 16'hF588;
defparam \Mux48~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N2
cycloneive_lcell_comb \Mux48~16 (
// Equation(s):
// \Mux48~16_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux48~13_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & (\Mux48~15_combout )))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux48~15_combout ),
	.datad(\Mux48~13_combout ),
	.cin(gnd),
	.combout(\Mux48~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~16 .lut_mask = 16'hBA98;
defparam \Mux48~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N25
dffeas \regs[3][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][15] .is_wysiwyg = "true";
defparam \regs[3][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N24
cycloneive_lcell_comb \Mux16~14 (
// Equation(s):
// \Mux16~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][15]~q ))) # (!dcifimemload_22 & (\regs[1][15]~q ))))

	.dataa(dcifimemload_22),
	.datab(\regs[1][15]~q ),
	.datac(\regs[3][15]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux16~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~14 .lut_mask = 16'hE400;
defparam \Mux16~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N16
cycloneive_lcell_comb \Mux16~15 (
// Equation(s):
// \Mux16~15_combout  = (\Mux16~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][15]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[2][15]~q ),
	.datad(\Mux16~14_combout ),
	.cin(gnd),
	.combout(\Mux16~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~15 .lut_mask = 16'hFF20;
defparam \Mux16~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N20
cycloneive_lcell_comb \Mux16~12 (
// Equation(s):
// \Mux16~12_combout  = (dcifimemload_21 & (((\regs[5][15]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][15]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][15]~q ),
	.datac(\regs[5][15]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux16~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~12 .lut_mask = 16'hAAE4;
defparam \Mux16~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N6
cycloneive_lcell_comb \Mux16~13 (
// Equation(s):
// \Mux16~13_combout  = (dcifimemload_22 & ((\Mux16~12_combout  & (\regs[7][15]~q )) # (!\Mux16~12_combout  & ((\regs[6][15]~q ))))) # (!dcifimemload_22 & (((\Mux16~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[7][15]~q ),
	.datac(\regs[6][15]~q ),
	.datad(\Mux16~12_combout ),
	.cin(gnd),
	.combout(\Mux16~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~13 .lut_mask = 16'hDDA0;
defparam \Mux16~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N18
cycloneive_lcell_comb \Mux16~16 (
// Equation(s):
// \Mux16~16_combout  = (dcifimemload_23 & (((dcifimemload_24) # (\Mux16~13_combout )))) # (!dcifimemload_23 & (\Mux16~15_combout  & (!dcifimemload_24)))

	.dataa(dcifimemload_23),
	.datab(\Mux16~15_combout ),
	.datac(dcifimemload_24),
	.datad(\Mux16~13_combout ),
	.cin(gnd),
	.combout(\Mux16~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~16 .lut_mask = 16'hAEA4;
defparam \Mux16~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N20
cycloneive_lcell_comb \Mux16~18 (
// Equation(s):
// \Mux16~18_combout  = (\Mux16~17_combout  & ((\regs[15][15]~q ) # ((!dcifimemload_22)))) # (!\Mux16~17_combout  & (((\regs[14][15]~q  & dcifimemload_22))))

	.dataa(\Mux16~17_combout ),
	.datab(\regs[15][15]~q ),
	.datac(\regs[14][15]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux16~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~18 .lut_mask = 16'hD8AA;
defparam \Mux16~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N9
dffeas \regs[10][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][15] .is_wysiwyg = "true";
defparam \regs[10][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N8
cycloneive_lcell_comb \Mux16~10 (
// Equation(s):
// \Mux16~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][15]~q ))) # (!dcifimemload_22 & (\regs[8][15]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][15]~q ),
	.datac(\regs[10][15]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~10 .lut_mask = 16'hFA44;
defparam \Mux16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N12
cycloneive_lcell_comb \Mux16~11 (
// Equation(s):
// \Mux16~11_combout  = (\Mux16~10_combout  & ((\regs[11][15]~q ) # ((!dcifimemload_21)))) # (!\Mux16~10_combout  & (((\regs[9][15]~q  & dcifimemload_21))))

	.dataa(\regs[11][15]~q ),
	.datab(\regs[9][15]~q ),
	.datac(\Mux16~10_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux16~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~11 .lut_mask = 16'hACF0;
defparam \Mux16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N4
cycloneive_lcell_comb \Mux16~19 (
// Equation(s):
// \Mux16~19_combout  = (dcifimemload_24 & ((\Mux16~16_combout  & (\Mux16~18_combout )) # (!\Mux16~16_combout  & ((\Mux16~11_combout ))))) # (!dcifimemload_24 & (\Mux16~16_combout ))

	.dataa(dcifimemload_24),
	.datab(\Mux16~16_combout ),
	.datac(\Mux16~18_combout ),
	.datad(\Mux16~11_combout ),
	.cin(gnd),
	.combout(\Mux16~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~19 .lut_mask = 16'hE6C4;
defparam \Mux16~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N14
cycloneive_lcell_comb \Mux16~8 (
// Equation(s):
// \Mux16~8_combout  = (\Mux16~7_combout  & (((\regs[31][15]~q ) # (!dcifimemload_24)))) # (!\Mux16~7_combout  & (\regs[27][15]~q  & ((dcifimemload_24))))

	.dataa(\Mux16~7_combout ),
	.datab(\regs[27][15]~q ),
	.datac(\regs[31][15]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~8 .lut_mask = 16'hE4AA;
defparam \Mux16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N3
dffeas \regs[24][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~32_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][15] .is_wysiwyg = "true";
defparam \regs[24][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N2
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (dcifimemload_24 & (((\regs[24][15]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[16][15]~q  & ((!dcifimemload_23))))

	.dataa(\regs[16][15]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[24][15]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hCCE2;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N2
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// \Mux16~5_combout  = (dcifimemload_23 & ((\Mux16~4_combout  & (\regs[28][15]~q )) # (!\Mux16~4_combout  & ((\regs[20][15]~q ))))) # (!dcifimemload_23 & (((\Mux16~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[28][15]~q ),
	.datac(\regs[20][15]~q ),
	.datad(\Mux16~4_combout ),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hDDA0;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N4
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (dcifimemload_22 & ((\Mux16~3_combout ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((\Mux16~5_combout  & !dcifimemload_21))))

	.dataa(\Mux16~3_combout ),
	.datab(dcifimemload_22),
	.datac(\Mux16~5_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hCCB8;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N4
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (dcifimemload_23 & (((\regs[21][15]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[17][15]~q  & ((!dcifimemload_24))))

	.dataa(\regs[17][15]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[21][15]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hCCE2;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N14
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (dcifimemload_24 & ((\Mux16~0_combout  & ((\regs[29][15]~q ))) # (!\Mux16~0_combout  & (\regs[25][15]~q )))) # (!dcifimemload_24 & (((\Mux16~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[25][15]~q ),
	.datac(\regs[29][15]~q ),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hF588;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N8
cycloneive_lcell_comb \Mux16~9 (
// Equation(s):
// \Mux16~9_combout  = (dcifimemload_21 & ((\Mux16~6_combout  & (\Mux16~8_combout )) # (!\Mux16~6_combout  & ((\Mux16~1_combout ))))) # (!dcifimemload_21 & (((\Mux16~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux16~8_combout ),
	.datac(\Mux16~6_combout ),
	.datad(\Mux16~1_combout ),
	.cin(gnd),
	.combout(\Mux16~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~9 .lut_mask = 16'hDAD0;
defparam \Mux16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N4
cycloneive_lcell_comb \regs~33 (
// Equation(s):
// \regs~33_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_14)) # (!cuifRegSel_0 & ((Mux173)))))

	.dataa(cuifRegSel_0),
	.datab(cuifRegSel_11),
	.datac(ramiframload_14),
	.datad(Mux171),
	.cin(gnd),
	.combout(\regs~33_combout ),
	.cout());
// synopsys translate_off
defparam \regs~33 .lut_mask = 16'h3120;
defparam \regs~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N10
cycloneive_lcell_comb \regs~34 (
// Equation(s):
// \regs~34_combout  = (!\Equal0~1_combout  & ((\regs~33_combout ) # ((\regs~64_combout  & \Add1~24_combout ))))

	.dataa(\regs~64_combout ),
	.datab(\regs~33_combout ),
	.datac(Add112),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\regs~34_combout ),
	.cout());
// synopsys translate_off
defparam \regs~34 .lut_mask = 16'h00EC;
defparam \regs~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N4
cycloneive_lcell_comb \regs[29][14]~feeder (
// Equation(s):
// \regs[29][14]~feeder_combout  = \regs~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~34_combout ),
	.cin(gnd),
	.combout(\regs[29][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][14]~feeder .lut_mask = 16'hFF00;
defparam \regs[29][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N5
dffeas \regs[29][14] (
	.clk(CLK),
	.d(\regs[29][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][14] .is_wysiwyg = "true";
defparam \regs[29][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N11
dffeas \regs[25][14] (
	.clk(CLK),
	.d(\regs~34_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][14] .is_wysiwyg = "true";
defparam \regs[25][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N20
cycloneive_lcell_comb \regs[21][14]~feeder (
// Equation(s):
// \regs[21][14]~feeder_combout  = \regs~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~34_combout ),
	.cin(gnd),
	.combout(\regs[21][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][14]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N21
dffeas \regs[21][14] (
	.clk(CLK),
	.d(\regs[21][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][14] .is_wysiwyg = "true";
defparam \regs[21][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N15
dffeas \regs[17][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][14] .is_wysiwyg = "true";
defparam \regs[17][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N14
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[21][14]~q )) # (!dcifimemload_18 & ((\regs[17][14]~q )))))

	.dataa(dcifimemload_19),
	.datab(\regs[21][14]~q ),
	.datac(\regs[17][14]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hEE50;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N12
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (\Mux49~0_combout  & ((\regs[29][14]~q ) # ((!dcifimemload_19)))) # (!\Mux49~0_combout  & (((\regs[25][14]~q  & dcifimemload_19))))

	.dataa(\regs[29][14]~q ),
	.datab(\regs[25][14]~q ),
	.datac(\Mux49~0_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hACF0;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N21
dffeas \regs[20][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][14] .is_wysiwyg = "true";
defparam \regs[20][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N1
dffeas \regs[28][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][14] .is_wysiwyg = "true";
defparam \regs[28][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N8
cycloneive_lcell_comb \regs[24][14]~feeder (
// Equation(s):
// \regs[24][14]~feeder_combout  = \regs~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~34_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[24][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][14]~feeder .lut_mask = 16'hF0F0;
defparam \regs[24][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N9
dffeas \regs[24][14] (
	.clk(CLK),
	.d(\regs[24][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][14] .is_wysiwyg = "true";
defparam \regs[24][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N7
dffeas \regs[16][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][14] .is_wysiwyg = "true";
defparam \regs[16][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N6
cycloneive_lcell_comb \Mux49~4 (
// Equation(s):
// \Mux49~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[24][14]~q )) # (!dcifimemload_19 & ((\regs[16][14]~q )))))

	.dataa(dcifimemload_18),
	.datab(\regs[24][14]~q ),
	.datac(\regs[16][14]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~4 .lut_mask = 16'hEE50;
defparam \Mux49~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N0
cycloneive_lcell_comb \Mux49~5 (
// Equation(s):
// \Mux49~5_combout  = (dcifimemload_18 & ((\Mux49~4_combout  & ((\regs[28][14]~q ))) # (!\Mux49~4_combout  & (\regs[20][14]~q )))) # (!dcifimemload_18 & (((\Mux49~4_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[20][14]~q ),
	.datac(\regs[28][14]~q ),
	.datad(\Mux49~4_combout ),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~5 .lut_mask = 16'hF588;
defparam \Mux49~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N23
dffeas \regs[30][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][14] .is_wysiwyg = "true";
defparam \regs[30][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N21
dffeas \regs[18][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][14] .is_wysiwyg = "true";
defparam \regs[18][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N20
cycloneive_lcell_comb \Mux49~2 (
// Equation(s):
// \Mux49~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[26][14]~q )) # (!dcifimemload_19 & ((\regs[18][14]~q )))))

	.dataa(\regs[26][14]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][14]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~2 .lut_mask = 16'hEE30;
defparam \Mux49~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N22
cycloneive_lcell_comb \Mux49~3 (
// Equation(s):
// \Mux49~3_combout  = (dcifimemload_18 & ((\Mux49~2_combout  & ((\regs[30][14]~q ))) # (!\Mux49~2_combout  & (\regs[22][14]~q )))) # (!dcifimemload_18 & (((\Mux49~2_combout ))))

	.dataa(\regs[22][14]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[30][14]~q ),
	.datad(\Mux49~2_combout ),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~3 .lut_mask = 16'hF388;
defparam \Mux49~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N30
cycloneive_lcell_comb \Mux49~6 (
// Equation(s):
// \Mux49~6_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux49~3_combout ))) # (!dcifimemload_17 & (\Mux49~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux49~5_combout ),
	.datac(dcifimemload_17),
	.datad(\Mux49~3_combout ),
	.cin(gnd),
	.combout(\Mux49~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~6 .lut_mask = 16'hF4A4;
defparam \Mux49~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N25
dffeas \regs[27][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][14] .is_wysiwyg = "true";
defparam \regs[27][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N15
dffeas \regs[31][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][14] .is_wysiwyg = "true";
defparam \regs[31][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N29
dffeas \regs[23][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][14] .is_wysiwyg = "true";
defparam \regs[23][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N19
dffeas \regs[19][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][14] .is_wysiwyg = "true";
defparam \regs[19][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N18
cycloneive_lcell_comb \Mux49~7 (
// Equation(s):
// \Mux49~7_combout  = (dcifimemload_18 & ((\regs[23][14]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[19][14]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[23][14]~q ),
	.datac(\regs[19][14]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux49~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~7 .lut_mask = 16'hAAD8;
defparam \Mux49~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N14
cycloneive_lcell_comb \Mux49~8 (
// Equation(s):
// \Mux49~8_combout  = (dcifimemload_19 & ((\Mux49~7_combout  & ((\regs[31][14]~q ))) # (!\Mux49~7_combout  & (\regs[27][14]~q )))) # (!dcifimemload_19 & (((\Mux49~7_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[27][14]~q ),
	.datac(\regs[31][14]~q ),
	.datad(\Mux49~7_combout ),
	.cin(gnd),
	.combout(\Mux49~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~8 .lut_mask = 16'hF588;
defparam \Mux49~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N11
dffeas \regs[9][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][14] .is_wysiwyg = "true";
defparam \regs[9][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N15
dffeas \regs[11][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][14] .is_wysiwyg = "true";
defparam \regs[11][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N31
dffeas \regs[10][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][14] .is_wysiwyg = "true";
defparam \regs[10][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N25
dffeas \regs[8][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][14] .is_wysiwyg = "true";
defparam \regs[8][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N24
cycloneive_lcell_comb \Mux49~10 (
// Equation(s):
// \Mux49~10_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][14]~q )) # (!dcifimemload_17 & ((\regs[8][14]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][14]~q ),
	.datac(\regs[8][14]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux49~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~10 .lut_mask = 16'hEE50;
defparam \Mux49~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N14
cycloneive_lcell_comb \Mux49~11 (
// Equation(s):
// \Mux49~11_combout  = (dcifimemload_16 & ((\Mux49~10_combout  & ((\regs[11][14]~q ))) # (!\Mux49~10_combout  & (\regs[9][14]~q )))) # (!dcifimemload_16 & (((\Mux49~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][14]~q ),
	.datac(\regs[11][14]~q ),
	.datad(\Mux49~10_combout ),
	.cin(gnd),
	.combout(\Mux49~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~11 .lut_mask = 16'hF588;
defparam \Mux49~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N10
cycloneive_lcell_comb \regs[15][14]~feeder (
// Equation(s):
// \regs[15][14]~feeder_combout  = \regs~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~34_combout ),
	.cin(gnd),
	.combout(\regs[15][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][14]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N11
dffeas \regs[15][14] (
	.clk(CLK),
	.d(\regs[15][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][14] .is_wysiwyg = "true";
defparam \regs[15][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N5
dffeas \regs[14][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][14] .is_wysiwyg = "true";
defparam \regs[14][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N16
cycloneive_lcell_comb \regs[12][14]~feeder (
// Equation(s):
// \regs[12][14]~feeder_combout  = \regs~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~34_combout ),
	.cin(gnd),
	.combout(\regs[12][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[12][14]~feeder .lut_mask = 16'hFF00;
defparam \regs[12][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N17
dffeas \regs[12][14] (
	.clk(CLK),
	.d(\regs[12][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][14] .is_wysiwyg = "true";
defparam \regs[12][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N22
cycloneive_lcell_comb \Mux49~17 (
// Equation(s):
// \Mux49~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][14]~q )) # (!dcifimemload_16 & ((\regs[12][14]~q )))))

	.dataa(\regs[13][14]~q ),
	.datab(\regs[12][14]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux49~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~17 .lut_mask = 16'hFA0C;
defparam \Mux49~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N16
cycloneive_lcell_comb \Mux49~18 (
// Equation(s):
// \Mux49~18_combout  = (dcifimemload_17 & ((\Mux49~17_combout  & (\regs[15][14]~q )) # (!\Mux49~17_combout  & ((\regs[14][14]~q ))))) # (!dcifimemload_17 & (((\Mux49~17_combout ))))

	.dataa(\regs[15][14]~q ),
	.datab(\regs[14][14]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux49~17_combout ),
	.cin(gnd),
	.combout(\Mux49~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~18 .lut_mask = 16'hAFC0;
defparam \Mux49~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N15
dffeas \regs[6][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][14] .is_wysiwyg = "true";
defparam \regs[6][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N21
dffeas \regs[7][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][14] .is_wysiwyg = "true";
defparam \regs[7][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N20
cycloneive_lcell_comb \Mux49~13 (
// Equation(s):
// \Mux49~13_combout  = (\Mux49~12_combout  & (((\regs[7][14]~q ) # (!dcifimemload_17)))) # (!\Mux49~12_combout  & (\regs[6][14]~q  & ((dcifimemload_17))))

	.dataa(\Mux49~12_combout ),
	.datab(\regs[6][14]~q ),
	.datac(\regs[7][14]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux49~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~13 .lut_mask = 16'hE4AA;
defparam \Mux49~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N5
dffeas \regs[2][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][14] .is_wysiwyg = "true";
defparam \regs[2][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N15
dffeas \regs[1][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][14] .is_wysiwyg = "true";
defparam \regs[1][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N13
dffeas \regs[3][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][14] .is_wysiwyg = "true";
defparam \regs[3][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N14
cycloneive_lcell_comb \Mux49~14 (
// Equation(s):
// \Mux49~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\regs[3][14]~q ))) # (!dcifimemload_17 & (\regs[1][14]~q ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[1][14]~q ),
	.datad(\regs[3][14]~q ),
	.cin(gnd),
	.combout(\Mux49~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~14 .lut_mask = 16'hA820;
defparam \Mux49~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N22
cycloneive_lcell_comb \Mux49~15 (
// Equation(s):
// \Mux49~15_combout  = (\Mux49~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][14]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][14]~q ),
	.datad(\Mux49~14_combout ),
	.cin(gnd),
	.combout(\Mux49~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~15 .lut_mask = 16'hFF40;
defparam \Mux49~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N10
cycloneive_lcell_comb \Mux49~16 (
// Equation(s):
// \Mux49~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & (\Mux49~13_combout )) # (!dcifimemload_18 & ((\Mux49~15_combout )))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux49~13_combout ),
	.datad(\Mux49~15_combout ),
	.cin(gnd),
	.combout(\Mux49~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~16 .lut_mask = 16'hD9C8;
defparam \Mux49~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N12
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[25][14]~q )) # (!dcifimemload_24 & ((\regs[17][14]~q )))))

	.dataa(\regs[25][14]~q ),
	.datab(\regs[17][14]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hFA0C;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N22
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (dcifimemload_23 & ((\Mux17~0_combout  & (\regs[29][14]~q )) # (!\Mux17~0_combout  & ((\regs[21][14]~q ))))) # (!dcifimemload_23 & (((\Mux17~0_combout ))))

	.dataa(\regs[29][14]~q ),
	.datab(\regs[21][14]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux17~0_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hAFC0;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N24
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// \Mux17~7_combout  = (dcifimemload_24 & (((\regs[27][14]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[19][14]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[19][14]~q ),
	.datac(\regs[27][14]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hAAE4;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N28
cycloneive_lcell_comb \Mux17~8 (
// Equation(s):
// \Mux17~8_combout  = (dcifimemload_23 & ((\Mux17~7_combout  & (\regs[31][14]~q )) # (!\Mux17~7_combout  & ((\regs[23][14]~q ))))) # (!dcifimemload_23 & (((\Mux17~7_combout ))))

	.dataa(\regs[31][14]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[23][14]~q ),
	.datad(\Mux17~7_combout ),
	.cin(gnd),
	.combout(\Mux17~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~8 .lut_mask = 16'hBBC0;
defparam \Mux17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N20
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[20][14]~q ))) # (!dcifimemload_23 & (\regs[16][14]~q ))))

	.dataa(\regs[16][14]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[20][14]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hFC22;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N30
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// \Mux17~5_combout  = (\Mux17~4_combout  & ((\regs[28][14]~q ) # ((!dcifimemload_24)))) # (!\Mux17~4_combout  & (((\regs[24][14]~q  & dcifimemload_24))))

	.dataa(\regs[28][14]~q ),
	.datab(\regs[24][14]~q ),
	.datac(\Mux17~4_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hACF0;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N24
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (dcifimemload_23 & ((\regs[22][14]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[18][14]~q  & !dcifimemload_24))))

	.dataa(\regs[22][14]~q ),
	.datab(\regs[18][14]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hF0AC;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N16
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (\Mux17~2_combout  & (((\regs[30][14]~q ) # (!dcifimemload_24)))) # (!\Mux17~2_combout  & (\regs[26][14]~q  & ((dcifimemload_24))))

	.dataa(\regs[26][14]~q ),
	.datab(\regs[30][14]~q ),
	.datac(\Mux17~2_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hCAF0;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N20
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// \Mux17~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux17~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux17~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux17~5_combout ),
	.datad(\Mux17~3_combout ),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'hBA98;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N26
cycloneive_lcell_comb \Mux17~9 (
// Equation(s):
// \Mux17~9_combout  = (dcifimemload_21 & ((\Mux17~6_combout  & ((\Mux17~8_combout ))) # (!\Mux17~6_combout  & (\Mux17~1_combout )))) # (!dcifimemload_21 & (((\Mux17~6_combout ))))

	.dataa(\Mux17~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux17~8_combout ),
	.datad(\Mux17~6_combout ),
	.cin(gnd),
	.combout(\Mux17~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~9 .lut_mask = 16'hF388;
defparam \Mux17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N12
cycloneive_lcell_comb \Mux17~14 (
// Equation(s):
// \Mux17~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][14]~q ))) # (!dcifimemload_22 & (\regs[1][14]~q ))))

	.dataa(\regs[1][14]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[3][14]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~14 .lut_mask = 16'hC088;
defparam \Mux17~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N4
cycloneive_lcell_comb \Mux17~15 (
// Equation(s):
// \Mux17~15_combout  = (\Mux17~14_combout ) # ((dcifimemload_22 & (\regs[2][14]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\regs[2][14]~q ),
	.datac(\Mux17~14_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux17~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~15 .lut_mask = 16'hF0F8;
defparam \Mux17~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \Mux17~12 (
// Equation(s):
// \Mux17~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][14]~q ))) # (!dcifimemload_22 & (\regs[8][14]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][14]~q ),
	.datac(\regs[10][14]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~12 .lut_mask = 16'hFA44;
defparam \Mux17~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N0
cycloneive_lcell_comb \Mux17~13 (
// Equation(s):
// \Mux17~13_combout  = (dcifimemload_21 & ((\Mux17~12_combout  & ((\regs[11][14]~q ))) # (!\Mux17~12_combout  & (\regs[9][14]~q )))) # (!dcifimemload_21 & (((\Mux17~12_combout ))))

	.dataa(\regs[9][14]~q ),
	.datab(\regs[11][14]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux17~12_combout ),
	.cin(gnd),
	.combout(\Mux17~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~13 .lut_mask = 16'hCFA0;
defparam \Mux17~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N18
cycloneive_lcell_comb \Mux17~16 (
// Equation(s):
// \Mux17~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux17~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & (\Mux17~15_combout )))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux17~15_combout ),
	.datad(\Mux17~13_combout ),
	.cin(gnd),
	.combout(\Mux17~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~16 .lut_mask = 16'hBA98;
defparam \Mux17~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N4
cycloneive_lcell_comb \Mux17~18 (
// Equation(s):
// \Mux17~18_combout  = (\Mux17~17_combout  & ((\regs[15][14]~q ) # ((!dcifimemload_22)))) # (!\Mux17~17_combout  & (((\regs[14][14]~q  & dcifimemload_22))))

	.dataa(\Mux17~17_combout ),
	.datab(\regs[15][14]~q ),
	.datac(\regs[14][14]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~18 .lut_mask = 16'hD8AA;
defparam \Mux17~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N7
dffeas \regs[4][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][14] .is_wysiwyg = "true";
defparam \regs[4][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N17
dffeas \regs[5][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~34_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][14] .is_wysiwyg = "true";
defparam \regs[5][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N16
cycloneive_lcell_comb \Mux17~10 (
// Equation(s):
// \Mux17~10_combout  = (dcifimemload_21 & (((\regs[5][14]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][14]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][14]~q ),
	.datac(\regs[5][14]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~10 .lut_mask = 16'hAAE4;
defparam \Mux17~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N14
cycloneive_lcell_comb \Mux17~11 (
// Equation(s):
// \Mux17~11_combout  = (\Mux17~10_combout  & ((\regs[7][14]~q ) # ((!dcifimemload_22)))) # (!\Mux17~10_combout  & (((\regs[6][14]~q  & dcifimemload_22))))

	.dataa(\regs[7][14]~q ),
	.datab(\Mux17~10_combout ),
	.datac(\regs[6][14]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~11 .lut_mask = 16'hB8CC;
defparam \Mux17~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N28
cycloneive_lcell_comb \Mux17~19 (
// Equation(s):
// \Mux17~19_combout  = (dcifimemload_23 & ((\Mux17~16_combout  & (\Mux17~18_combout )) # (!\Mux17~16_combout  & ((\Mux17~11_combout ))))) # (!dcifimemload_23 & (\Mux17~16_combout ))

	.dataa(dcifimemload_23),
	.datab(\Mux17~16_combout ),
	.datac(\Mux17~18_combout ),
	.datad(\Mux17~11_combout ),
	.cin(gnd),
	.combout(\Mux17~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~19 .lut_mask = 16'hE6C4;
defparam \Mux17~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N10
cycloneive_lcell_comb \regs~35 (
// Equation(s):
// \regs~35_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_13)) # (!cuifRegSel_0 & ((Mux183)))))

	.dataa(cuifRegSel_0),
	.datab(cuifRegSel_11),
	.datac(ramiframload_13),
	.datad(Mux181),
	.cin(gnd),
	.combout(\regs~35_combout ),
	.cout());
// synopsys translate_off
defparam \regs~35 .lut_mask = 16'h3120;
defparam \regs~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N24
cycloneive_lcell_comb \regs~36 (
// Equation(s):
// \regs~36_combout  = (!\Equal0~1_combout  & ((\regs~35_combout ) # ((\regs~64_combout  & \Add1~22_combout ))))

	.dataa(\regs~64_combout ),
	.datab(Add111),
	.datac(\Equal0~1_combout ),
	.datad(\regs~35_combout ),
	.cin(gnd),
	.combout(\regs~36_combout ),
	.cout());
// synopsys translate_off
defparam \regs~36 .lut_mask = 16'h0F08;
defparam \regs~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N15
dffeas \regs[23][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][13] .is_wysiwyg = "true";
defparam \regs[23][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N3
dffeas \regs[31][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][13] .is_wysiwyg = "true";
defparam \regs[31][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N0
cycloneive_lcell_comb \regs[19][13]~feeder (
// Equation(s):
// \regs[19][13]~feeder_combout  = \regs~36_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~36_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[19][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][13]~feeder .lut_mask = 16'hF0F0;
defparam \regs[19][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N1
dffeas \regs[19][13] (
	.clk(CLK),
	.d(\regs[19][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][13] .is_wysiwyg = "true";
defparam \regs[19][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N16
cycloneive_lcell_comb \Mux50~7 (
// Equation(s):
// \Mux50~7_combout  = (dcifimemload_19 & ((\regs[27][13]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\regs[19][13]~q  & !dcifimemload_18))))

	.dataa(\regs[27][13]~q ),
	.datab(\regs[19][13]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux50~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~7 .lut_mask = 16'hF0AC;
defparam \Mux50~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N2
cycloneive_lcell_comb \Mux50~8 (
// Equation(s):
// \Mux50~8_combout  = (dcifimemload_18 & ((\Mux50~7_combout  & ((\regs[31][13]~q ))) # (!\Mux50~7_combout  & (\regs[23][13]~q )))) # (!dcifimemload_18 & (((\Mux50~7_combout ))))

	.dataa(\regs[23][13]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[31][13]~q ),
	.datad(\Mux50~7_combout ),
	.cin(gnd),
	.combout(\Mux50~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~8 .lut_mask = 16'hF388;
defparam \Mux50~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N5
dffeas \regs[18][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][13] .is_wysiwyg = "true";
defparam \regs[18][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N4
cycloneive_lcell_comb \Mux50~2 (
// Equation(s):
// \Mux50~2_combout  = (dcifimemload_18 & ((\regs[22][13]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[18][13]~q  & !dcifimemload_19))))

	.dataa(\regs[22][13]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][13]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~2 .lut_mask = 16'hCCB8;
defparam \Mux50~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N31
dffeas \regs[30][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][13] .is_wysiwyg = "true";
defparam \regs[30][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N30
cycloneive_lcell_comb \Mux50~3 (
// Equation(s):
// \Mux50~3_combout  = (\Mux50~2_combout  & (((\regs[30][13]~q ) # (!dcifimemload_19)))) # (!\Mux50~2_combout  & (\regs[26][13]~q  & ((dcifimemload_19))))

	.dataa(\regs[26][13]~q ),
	.datab(\Mux50~2_combout ),
	.datac(\regs[30][13]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~3 .lut_mask = 16'hE2CC;
defparam \Mux50~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N13
dffeas \regs[24][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][13] .is_wysiwyg = "true";
defparam \regs[24][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N23
dffeas \regs[28][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][13] .is_wysiwyg = "true";
defparam \regs[28][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N1
dffeas \regs[16][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][13] .is_wysiwyg = "true";
defparam \regs[16][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N0
cycloneive_lcell_comb \Mux50~4 (
// Equation(s):
// \Mux50~4_combout  = (dcifimemload_18 & ((\regs[20][13]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[16][13]~q  & !dcifimemload_19))))

	.dataa(\regs[20][13]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[16][13]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux50~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~4 .lut_mask = 16'hCCB8;
defparam \Mux50~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N22
cycloneive_lcell_comb \Mux50~5 (
// Equation(s):
// \Mux50~5_combout  = (dcifimemload_19 & ((\Mux50~4_combout  & ((\regs[28][13]~q ))) # (!\Mux50~4_combout  & (\regs[24][13]~q )))) # (!dcifimemload_19 & (((\Mux50~4_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[24][13]~q ),
	.datac(\regs[28][13]~q ),
	.datad(\Mux50~4_combout ),
	.cin(gnd),
	.combout(\Mux50~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~5 .lut_mask = 16'hF588;
defparam \Mux50~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N8
cycloneive_lcell_comb \Mux50~6 (
// Equation(s):
// \Mux50~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux50~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & ((\Mux50~5_combout ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux50~3_combout ),
	.datad(\Mux50~5_combout ),
	.cin(gnd),
	.combout(\Mux50~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~6 .lut_mask = 16'hB9A8;
defparam \Mux50~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N25
dffeas \regs[21][13] (
	.clk(CLK),
	.d(\regs~36_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][13] .is_wysiwyg = "true";
defparam \regs[21][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N8
cycloneive_lcell_comb \regs[29][13]~feeder (
// Equation(s):
// \regs[29][13]~feeder_combout  = \regs~36_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~36_combout ),
	.cin(gnd),
	.combout(\regs[29][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[29][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N9
dffeas \regs[29][13] (
	.clk(CLK),
	.d(\regs[29][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][13] .is_wysiwyg = "true";
defparam \regs[29][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N19
dffeas \regs[25][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][13] .is_wysiwyg = "true";
defparam \regs[25][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N21
dffeas \regs[17][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][13] .is_wysiwyg = "true";
defparam \regs[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N18
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[25][13]~q )) # (!dcifimemload_19 & ((\regs[17][13]~q )))))

	.dataa(dcifimemload_18),
	.datab(\regs[25][13]~q ),
	.datac(\regs[17][13]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hEE50;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N30
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (dcifimemload_18 & ((\Mux50~0_combout  & ((\regs[29][13]~q ))) # (!\Mux50~0_combout  & (\regs[21][13]~q )))) # (!dcifimemload_18 & (((\Mux50~0_combout ))))

	.dataa(\regs[21][13]~q ),
	.datab(\regs[29][13]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux50~0_combout ),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hCFA0;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N12
cycloneive_lcell_comb \regs[15][13]~feeder (
// Equation(s):
// \regs[15][13]~feeder_combout  = \regs~36_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~36_combout ),
	.cin(gnd),
	.combout(\regs[15][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N13
dffeas \regs[15][13] (
	.clk(CLK),
	.d(\regs[15][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][13] .is_wysiwyg = "true";
defparam \regs[15][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N9
dffeas \regs[14][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][13] .is_wysiwyg = "true";
defparam \regs[14][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N7
dffeas \regs[13][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][13] .is_wysiwyg = "true";
defparam \regs[13][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N6
cycloneive_lcell_comb \Mux50~17 (
// Equation(s):
// \Mux50~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\regs[13][13]~q ))) # (!dcifimemload_16 & (\regs[12][13]~q ))))

	.dataa(\regs[12][13]~q ),
	.datab(\regs[13][13]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux50~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~17 .lut_mask = 16'hFC0A;
defparam \Mux50~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N22
cycloneive_lcell_comb \Mux50~18 (
// Equation(s):
// \Mux50~18_combout  = (dcifimemload_17 & ((\Mux50~17_combout  & (\regs[15][13]~q )) # (!\Mux50~17_combout  & ((\regs[14][13]~q ))))) # (!dcifimemload_17 & (((\Mux50~17_combout ))))

	.dataa(\regs[15][13]~q ),
	.datab(\regs[14][13]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux50~17_combout ),
	.cin(gnd),
	.combout(\Mux50~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~18 .lut_mask = 16'hAFC0;
defparam \Mux50~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N23
dffeas \regs[6][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][13] .is_wysiwyg = "true";
defparam \regs[6][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N9
dffeas \regs[7][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][13] .is_wysiwyg = "true";
defparam \regs[7][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N13
dffeas \regs[5][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][13] .is_wysiwyg = "true";
defparam \regs[5][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N23
dffeas \regs[4][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][13] .is_wysiwyg = "true";
defparam \regs[4][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N22
cycloneive_lcell_comb \Mux50~10 (
// Equation(s):
// \Mux50~10_combout  = (dcifimemload_16 & ((\regs[5][13]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][13]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[5][13]~q ),
	.datac(\regs[4][13]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux50~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~10 .lut_mask = 16'hAAD8;
defparam \Mux50~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N10
cycloneive_lcell_comb \Mux50~11 (
// Equation(s):
// \Mux50~11_combout  = (dcifimemload_17 & ((\Mux50~10_combout  & ((\regs[7][13]~q ))) # (!\Mux50~10_combout  & (\regs[6][13]~q )))) # (!dcifimemload_17 & (((\Mux50~10_combout ))))

	.dataa(\regs[6][13]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[7][13]~q ),
	.datad(\Mux50~10_combout ),
	.cin(gnd),
	.combout(\Mux50~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~11 .lut_mask = 16'hF388;
defparam \Mux50~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N4
cycloneive_lcell_comb \regs[9][13]~feeder (
// Equation(s):
// \regs[9][13]~feeder_combout  = \regs~36_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~36_combout ),
	.cin(gnd),
	.combout(\regs[9][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N5
dffeas \regs[9][13] (
	.clk(CLK),
	.d(\regs[9][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][13] .is_wysiwyg = "true";
defparam \regs[9][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N27
dffeas \regs[11][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][13] .is_wysiwyg = "true";
defparam \regs[11][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N31
dffeas \regs[10][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][13] .is_wysiwyg = "true";
defparam \regs[10][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N13
dffeas \regs[8][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][13] .is_wysiwyg = "true";
defparam \regs[8][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N12
cycloneive_lcell_comb \Mux50~12 (
// Equation(s):
// \Mux50~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][13]~q )) # (!dcifimemload_17 & ((\regs[8][13]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][13]~q ),
	.datac(\regs[8][13]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux50~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~12 .lut_mask = 16'hEE50;
defparam \Mux50~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N26
cycloneive_lcell_comb \Mux50~13 (
// Equation(s):
// \Mux50~13_combout  = (dcifimemload_16 & ((\Mux50~12_combout  & ((\regs[11][13]~q ))) # (!\Mux50~12_combout  & (\regs[9][13]~q )))) # (!dcifimemload_16 & (((\Mux50~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][13]~q ),
	.datac(\regs[11][13]~q ),
	.datad(\Mux50~12_combout ),
	.cin(gnd),
	.combout(\Mux50~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~13 .lut_mask = 16'hF588;
defparam \Mux50~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N31
dffeas \regs[2][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][13] .is_wysiwyg = "true";
defparam \regs[2][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N13
dffeas \regs[1][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][13] .is_wysiwyg = "true";
defparam \regs[1][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N12
cycloneive_lcell_comb \Mux50~14 (
// Equation(s):
// \Mux50~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][13]~q )) # (!dcifimemload_17 & ((\regs[1][13]~q )))))

	.dataa(\regs[3][13]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][13]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux50~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~14 .lut_mask = 16'h88C0;
defparam \Mux50~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N30
cycloneive_lcell_comb \Mux50~15 (
// Equation(s):
// \Mux50~15_combout  = (\Mux50~14_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][13]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[2][13]~q ),
	.datad(\Mux50~14_combout ),
	.cin(gnd),
	.combout(\Mux50~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~15 .lut_mask = 16'hFF20;
defparam \Mux50~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N20
cycloneive_lcell_comb \Mux50~16 (
// Equation(s):
// \Mux50~16_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux50~13_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & ((\Mux50~15_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux50~13_combout ),
	.datad(\Mux50~15_combout ),
	.cin(gnd),
	.combout(\Mux50~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~16 .lut_mask = 16'hB9A8;
defparam \Mux50~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N20
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[21][13]~q )) # (!dcifimemload_23 & ((\regs[17][13]~q )))))

	.dataa(\regs[21][13]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[17][13]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hEE30;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N18
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (dcifimemload_24 & ((\Mux18~0_combout  & (\regs[29][13]~q )) # (!\Mux18~0_combout  & ((\regs[25][13]~q ))))) # (!dcifimemload_24 & (((\Mux18~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[29][13]~q ),
	.datac(\regs[25][13]~q ),
	.datad(\Mux18~0_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hDDA0;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N19
dffeas \regs[20][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][13] .is_wysiwyg = "true";
defparam \regs[20][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N12
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (dcifimemload_24 & (((\regs[24][13]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[16][13]~q  & ((!dcifimemload_23))))

	.dataa(\regs[16][13]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[24][13]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hCCE2;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N18
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (dcifimemload_23 & ((\Mux18~4_combout  & (\regs[28][13]~q )) # (!\Mux18~4_combout  & ((\regs[20][13]~q ))))) # (!dcifimemload_23 & (((\Mux18~4_combout ))))

	.dataa(\regs[28][13]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[20][13]~q ),
	.datad(\Mux18~4_combout ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hBBC0;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N25
dffeas \regs[22][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][13] .is_wysiwyg = "true";
defparam \regs[22][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N29
dffeas \regs[26][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][13] .is_wysiwyg = "true";
defparam \regs[26][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N28
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\regs[26][13]~q ))) # (!dcifimemload_24 & (\regs[18][13]~q ))))

	.dataa(dcifimemload_23),
	.datab(\regs[18][13]~q ),
	.datac(\regs[26][13]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hFA44;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N24
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (dcifimemload_23 & ((\Mux18~2_combout  & (\regs[30][13]~q )) # (!\Mux18~2_combout  & ((\regs[22][13]~q ))))) # (!dcifimemload_23 & (((\Mux18~2_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[30][13]~q ),
	.datac(\regs[22][13]~q ),
	.datad(\Mux18~2_combout ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hDDA0;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N4
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux18~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux18~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux18~5_combout ),
	.datad(\Mux18~3_combout ),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hBA98;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N27
dffeas \regs[27][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~36_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][13] .is_wysiwyg = "true";
defparam \regs[27][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N14
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (dcifimemload_23 & (((\regs[23][13]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[19][13]~q  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[19][13]~q ),
	.datac(\regs[23][13]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hAAE4;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N26
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// \Mux18~8_combout  = (dcifimemload_24 & ((\Mux18~7_combout  & (\regs[31][13]~q )) # (!\Mux18~7_combout  & ((\regs[27][13]~q ))))) # (!dcifimemload_24 & (((\Mux18~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[31][13]~q ),
	.datac(\regs[27][13]~q ),
	.datad(\Mux18~7_combout ),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hDDA0;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N26
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// \Mux18~9_combout  = (dcifimemload_21 & ((\Mux18~6_combout  & ((\Mux18~8_combout ))) # (!\Mux18~6_combout  & (\Mux18~1_combout )))) # (!dcifimemload_21 & (((\Mux18~6_combout ))))

	.dataa(\Mux18~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux18~6_combout ),
	.datad(\Mux18~8_combout ),
	.cin(gnd),
	.combout(\Mux18~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'hF838;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N28
cycloneive_lcell_comb \regs[12][13]~feeder (
// Equation(s):
// \regs[12][13]~feeder_combout  = \regs~36_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~36_combout ),
	.cin(gnd),
	.combout(\regs[12][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[12][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[12][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N29
dffeas \regs[12][13] (
	.clk(CLK),
	.d(\regs[12][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][13] .is_wysiwyg = "true";
defparam \regs[12][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N6
cycloneive_lcell_comb \Mux18~17 (
// Equation(s):
// \Mux18~17_combout  = (dcifimemload_21 & (((\regs[13][13]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][13]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][13]~q ),
	.datac(\regs[13][13]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux18~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~17 .lut_mask = 16'hAAE4;
defparam \Mux18~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N8
cycloneive_lcell_comb \Mux18~18 (
// Equation(s):
// \Mux18~18_combout  = (dcifimemload_22 & ((\Mux18~17_combout  & (\regs[15][13]~q )) # (!\Mux18~17_combout  & ((\regs[14][13]~q ))))) # (!dcifimemload_22 & (((\Mux18~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][13]~q ),
	.datac(\regs[14][13]~q ),
	.datad(\Mux18~17_combout ),
	.cin(gnd),
	.combout(\Mux18~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~18 .lut_mask = 16'hDDA0;
defparam \Mux18~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N30
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// \Mux18~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][13]~q ))) # (!dcifimemload_22 & (\regs[8][13]~q ))))

	.dataa(\regs[8][13]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[10][13]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hFC22;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N18
cycloneive_lcell_comb \Mux18~11 (
// Equation(s):
// \Mux18~11_combout  = (dcifimemload_21 & ((\Mux18~10_combout  & (\regs[11][13]~q )) # (!\Mux18~10_combout  & ((\regs[9][13]~q ))))) # (!dcifimemload_21 & (((\Mux18~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\regs[11][13]~q ),
	.datac(\regs[9][13]~q ),
	.datad(\Mux18~10_combout ),
	.cin(gnd),
	.combout(\Mux18~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~11 .lut_mask = 16'hDDA0;
defparam \Mux18~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N12
cycloneive_lcell_comb \Mux18~12 (
// Equation(s):
// \Mux18~12_combout  = (dcifimemload_21 & (((\regs[5][13]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][13]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][13]~q ),
	.datac(\regs[5][13]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux18~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~12 .lut_mask = 16'hAAE4;
defparam \Mux18~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N22
cycloneive_lcell_comb \Mux18~13 (
// Equation(s):
// \Mux18~13_combout  = (dcifimemload_22 & ((\Mux18~12_combout  & (\regs[7][13]~q )) # (!\Mux18~12_combout  & ((\regs[6][13]~q ))))) # (!dcifimemload_22 & (((\Mux18~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[7][13]~q ),
	.datac(\regs[6][13]~q ),
	.datad(\Mux18~12_combout ),
	.cin(gnd),
	.combout(\Mux18~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~13 .lut_mask = 16'hDDA0;
defparam \Mux18~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N20
cycloneive_lcell_comb \Mux18~14 (
// Equation(s):
// \Mux18~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\regs[3][13]~q )) # (!dcifimemload_22 & ((\regs[1][13]~q )))))

	.dataa(\regs[3][13]~q ),
	.datab(\regs[1][13]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux18~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~14 .lut_mask = 16'hA0C0;
defparam \Mux18~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N24
cycloneive_lcell_comb \Mux18~15 (
// Equation(s):
// \Mux18~15_combout  = (\Mux18~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][13]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[2][13]~q ),
	.datad(\Mux18~14_combout ),
	.cin(gnd),
	.combout(\Mux18~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~15 .lut_mask = 16'hFF20;
defparam \Mux18~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N18
cycloneive_lcell_comb \Mux18~16 (
// Equation(s):
// \Mux18~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux18~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & ((\Mux18~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux18~13_combout ),
	.datad(\Mux18~15_combout ),
	.cin(gnd),
	.combout(\Mux18~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~16 .lut_mask = 16'hB9A8;
defparam \Mux18~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N28
cycloneive_lcell_comb \Mux18~19 (
// Equation(s):
// \Mux18~19_combout  = (dcifimemload_24 & ((\Mux18~16_combout  & (\Mux18~18_combout )) # (!\Mux18~16_combout  & ((\Mux18~11_combout ))))) # (!dcifimemload_24 & (((\Mux18~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux18~18_combout ),
	.datac(\Mux18~11_combout ),
	.datad(\Mux18~16_combout ),
	.cin(gnd),
	.combout(\Mux18~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~19 .lut_mask = 16'hDDA0;
defparam \Mux18~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N30
cycloneive_lcell_comb \regs~37 (
// Equation(s):
// \regs~37_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_12)) # (!cuifRegSel_0 & ((Mux193)))))

	.dataa(ramiframload_12),
	.datab(cuifRegSel_11),
	.datac(Mux191),
	.datad(cuifRegSel_0),
	.cin(gnd),
	.combout(\regs~37_combout ),
	.cout());
// synopsys translate_off
defparam \regs~37 .lut_mask = 16'h2230;
defparam \regs~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N22
cycloneive_lcell_comb \regs~38 (
// Equation(s):
// \regs~38_combout  = (!\Equal0~1_combout  & ((\regs~37_combout ) # ((\regs~64_combout  & \Add1~20_combout ))))

	.dataa(\regs~64_combout ),
	.datab(Add110),
	.datac(\regs~37_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\regs~38_combout ),
	.cout());
// synopsys translate_off
defparam \regs~38 .lut_mask = 16'h00F8;
defparam \regs~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N30
cycloneive_lcell_comb \regs[31][12]~feeder (
// Equation(s):
// \regs[31][12]~feeder_combout  = \regs~38_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~38_combout ),
	.cin(gnd),
	.combout(\regs[31][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][12]~feeder .lut_mask = 16'hFF00;
defparam \regs[31][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N31
dffeas \regs[31][12] (
	.clk(CLK),
	.d(\regs[31][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][12] .is_wysiwyg = "true";
defparam \regs[31][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N5
dffeas \regs[27][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][12] .is_wysiwyg = "true";
defparam \regs[27][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N21
dffeas \regs[19][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][12] .is_wysiwyg = "true";
defparam \regs[19][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N27
dffeas \regs[23][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][12] .is_wysiwyg = "true";
defparam \regs[23][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N20
cycloneive_lcell_comb \Mux51~7 (
// Equation(s):
// \Mux51~7_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\regs[23][12]~q )))) # (!dcifimemload_18 & (!dcifimemload_19 & (\regs[19][12]~q )))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\regs[19][12]~q ),
	.datad(\regs[23][12]~q ),
	.cin(gnd),
	.combout(\Mux51~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~7 .lut_mask = 16'hBA98;
defparam \Mux51~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N6
cycloneive_lcell_comb \Mux51~8 (
// Equation(s):
// \Mux51~8_combout  = (dcifimemload_19 & ((\Mux51~7_combout  & (\regs[31][12]~q )) # (!\Mux51~7_combout  & ((\regs[27][12]~q ))))) # (!dcifimemload_19 & (((\Mux51~7_combout ))))

	.dataa(\regs[31][12]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[27][12]~q ),
	.datad(\Mux51~7_combout ),
	.cin(gnd),
	.combout(\Mux51~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~8 .lut_mask = 16'hBBC0;
defparam \Mux51~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N21
dffeas \regs[21][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][12] .is_wysiwyg = "true";
defparam \regs[21][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N23
dffeas \regs[17][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][12] .is_wysiwyg = "true";
defparam \regs[17][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N22
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (dcifimemload_18 & ((\regs[21][12]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[17][12]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[21][12]~q ),
	.datac(\regs[17][12]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hAAD8;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N23
dffeas \regs[25][12] (
	.clk(CLK),
	.d(\regs~38_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][12] .is_wysiwyg = "true";
defparam \regs[25][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N13
dffeas \regs[29][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][12] .is_wysiwyg = "true";
defparam \regs[29][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N12
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (\Mux51~0_combout  & (((\regs[29][12]~q ) # (!dcifimemload_19)))) # (!\Mux51~0_combout  & (\regs[25][12]~q  & ((dcifimemload_19))))

	.dataa(\Mux51~0_combout ),
	.datab(\regs[25][12]~q ),
	.datac(\regs[29][12]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hE4AA;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N31
dffeas \regs[20][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][12] .is_wysiwyg = "true";
defparam \regs[20][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N3
dffeas \regs[28][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][12] .is_wysiwyg = "true";
defparam \regs[28][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N25
dffeas \regs[16][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][12] .is_wysiwyg = "true";
defparam \regs[16][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N24
cycloneive_lcell_comb \Mux51~4 (
// Equation(s):
// \Mux51~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[24][12]~q )) # (!dcifimemload_19 & ((\regs[16][12]~q )))))

	.dataa(\regs[24][12]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[16][12]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux51~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~4 .lut_mask = 16'hEE30;
defparam \Mux51~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N2
cycloneive_lcell_comb \Mux51~5 (
// Equation(s):
// \Mux51~5_combout  = (dcifimemload_18 & ((\Mux51~4_combout  & ((\regs[28][12]~q ))) # (!\Mux51~4_combout  & (\regs[20][12]~q )))) # (!dcifimemload_18 & (((\Mux51~4_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[20][12]~q ),
	.datac(\regs[28][12]~q ),
	.datad(\Mux51~4_combout ),
	.cin(gnd),
	.combout(\Mux51~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~5 .lut_mask = 16'hF588;
defparam \Mux51~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N15
dffeas \regs[30][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][12] .is_wysiwyg = "true";
defparam \regs[30][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N9
dffeas \regs[18][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][12] .is_wysiwyg = "true";
defparam \regs[18][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N8
cycloneive_lcell_comb \Mux51~2 (
// Equation(s):
// \Mux51~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[26][12]~q )) # (!dcifimemload_19 & ((\regs[18][12]~q )))))

	.dataa(\regs[26][12]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][12]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux51~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~2 .lut_mask = 16'hEE30;
defparam \Mux51~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N14
cycloneive_lcell_comb \Mux51~3 (
// Equation(s):
// \Mux51~3_combout  = (dcifimemload_18 & ((\Mux51~2_combout  & ((\regs[30][12]~q ))) # (!\Mux51~2_combout  & (\regs[22][12]~q )))) # (!dcifimemload_18 & (((\Mux51~2_combout ))))

	.dataa(\regs[22][12]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[30][12]~q ),
	.datad(\Mux51~2_combout ),
	.cin(gnd),
	.combout(\Mux51~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~3 .lut_mask = 16'hF388;
defparam \Mux51~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N16
cycloneive_lcell_comb \Mux51~6 (
// Equation(s):
// \Mux51~6_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux51~3_combout ))) # (!dcifimemload_17 & (\Mux51~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux51~5_combout ),
	.datac(dcifimemload_17),
	.datad(\Mux51~3_combout ),
	.cin(gnd),
	.combout(\Mux51~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~6 .lut_mask = 16'hF4A4;
defparam \Mux51~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N5
dffeas \regs[8][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][12] .is_wysiwyg = "true";
defparam \regs[8][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N13
dffeas \regs[10][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][12] .is_wysiwyg = "true";
defparam \regs[10][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N4
cycloneive_lcell_comb \Mux51~10 (
// Equation(s):
// \Mux51~10_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\regs[10][12]~q ))) # (!dcifimemload_17 & (\regs[8][12]~q ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[8][12]~q ),
	.datad(\regs[10][12]~q ),
	.cin(gnd),
	.combout(\Mux51~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~10 .lut_mask = 16'hDC98;
defparam \Mux51~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N19
dffeas \regs[11][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][12] .is_wysiwyg = "true";
defparam \regs[11][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N7
dffeas \regs[9][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][12] .is_wysiwyg = "true";
defparam \regs[9][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N18
cycloneive_lcell_comb \Mux51~11 (
// Equation(s):
// \Mux51~11_combout  = (dcifimemload_16 & ((\Mux51~10_combout  & (\regs[11][12]~q )) # (!\Mux51~10_combout  & ((\regs[9][12]~q ))))) # (!dcifimemload_16 & (\Mux51~10_combout ))

	.dataa(dcifimemload_16),
	.datab(\Mux51~10_combout ),
	.datac(\regs[11][12]~q ),
	.datad(\regs[9][12]~q ),
	.cin(gnd),
	.combout(\Mux51~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~11 .lut_mask = 16'hE6C4;
defparam \Mux51~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N16
cycloneive_lcell_comb \regs[14][12]~feeder (
// Equation(s):
// \regs[14][12]~feeder_combout  = \regs~38_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~38_combout ),
	.cin(gnd),
	.combout(\regs[14][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][12]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y44_N17
dffeas \regs[14][12] (
	.clk(CLK),
	.d(\regs[14][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][12] .is_wysiwyg = "true";
defparam \regs[14][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y44_N3
dffeas \regs[15][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][12] .is_wysiwyg = "true";
defparam \regs[15][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N13
dffeas \regs[13][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][12] .is_wysiwyg = "true";
defparam \regs[13][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N27
dffeas \regs[12][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][12] .is_wysiwyg = "true";
defparam \regs[12][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N26
cycloneive_lcell_comb \Mux51~17 (
// Equation(s):
// \Mux51~17_combout  = (dcifimemload_16 & ((\regs[13][12]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[12][12]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[13][12]~q ),
	.datac(\regs[12][12]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux51~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~17 .lut_mask = 16'hAAD8;
defparam \Mux51~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N2
cycloneive_lcell_comb \Mux51~18 (
// Equation(s):
// \Mux51~18_combout  = (dcifimemload_17 & ((\Mux51~17_combout  & ((\regs[15][12]~q ))) # (!\Mux51~17_combout  & (\regs[14][12]~q )))) # (!dcifimemload_17 & (((\Mux51~17_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[14][12]~q ),
	.datac(\regs[15][12]~q ),
	.datad(\Mux51~17_combout ),
	.cin(gnd),
	.combout(\Mux51~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~18 .lut_mask = 16'hF588;
defparam \Mux51~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N31
dffeas \regs[6][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][12] .is_wysiwyg = "true";
defparam \regs[6][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N11
dffeas \regs[7][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][12] .is_wysiwyg = "true";
defparam \regs[7][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N1
dffeas \regs[4][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][12] .is_wysiwyg = "true";
defparam \regs[4][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N0
cycloneive_lcell_comb \Mux51~12 (
// Equation(s):
// \Mux51~12_combout  = (dcifimemload_16 & ((\regs[5][12]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][12]~q  & !dcifimemload_17))))

	.dataa(\regs[5][12]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][12]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux51~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~12 .lut_mask = 16'hCCB8;
defparam \Mux51~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N10
cycloneive_lcell_comb \Mux51~13 (
// Equation(s):
// \Mux51~13_combout  = (dcifimemload_17 & ((\Mux51~12_combout  & ((\regs[7][12]~q ))) # (!\Mux51~12_combout  & (\regs[6][12]~q )))) # (!dcifimemload_17 & (((\Mux51~12_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][12]~q ),
	.datac(\regs[7][12]~q ),
	.datad(\Mux51~12_combout ),
	.cin(gnd),
	.combout(\Mux51~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~13 .lut_mask = 16'hF588;
defparam \Mux51~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y32_N23
dffeas \regs[2][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][12] .is_wysiwyg = "true";
defparam \regs[2][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N21
dffeas \regs[1][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][12] .is_wysiwyg = "true";
defparam \regs[1][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N20
cycloneive_lcell_comb \Mux51~14 (
// Equation(s):
// \Mux51~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][12]~q )) # (!dcifimemload_17 & ((\regs[1][12]~q )))))

	.dataa(\regs[3][12]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][12]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux51~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~14 .lut_mask = 16'h88C0;
defparam \Mux51~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N22
cycloneive_lcell_comb \Mux51~15 (
// Equation(s):
// \Mux51~15_combout  = (\Mux51~14_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][12]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[2][12]~q ),
	.datad(\Mux51~14_combout ),
	.cin(gnd),
	.combout(\Mux51~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~15 .lut_mask = 16'hFF20;
defparam \Mux51~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N24
cycloneive_lcell_comb \Mux51~16 (
// Equation(s):
// \Mux51~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & (\Mux51~13_combout )) # (!dcifimemload_18 & ((\Mux51~15_combout )))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux51~13_combout ),
	.datad(\Mux51~15_combout ),
	.cin(gnd),
	.combout(\Mux51~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~16 .lut_mask = 16'hD9C8;
defparam \Mux51~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N16
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (\Mux19~0_combout  & (((\regs[29][12]~q ) # (!dcifimemload_23)))) # (!\Mux19~0_combout  & (\regs[21][12]~q  & ((dcifimemload_23))))

	.dataa(\Mux19~0_combout ),
	.datab(\regs[21][12]~q ),
	.datac(\regs[29][12]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hE4AA;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N0
cycloneive_lcell_comb \regs[26][12]~feeder (
// Equation(s):
// \regs[26][12]~feeder_combout  = \regs~38_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~38_combout ),
	.cin(gnd),
	.combout(\regs[26][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][12]~feeder .lut_mask = 16'hFF00;
defparam \regs[26][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N1
dffeas \regs[26][12] (
	.clk(CLK),
	.d(\regs[26][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][12] .is_wysiwyg = "true";
defparam \regs[26][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N31
dffeas \regs[22][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][12] .is_wysiwyg = "true";
defparam \regs[22][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N30
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (dcifimemload_23 & (((\regs[22][12]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[18][12]~q  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[18][12]~q ),
	.datac(\regs[22][12]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hAAE4;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N28
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (\Mux19~2_combout  & ((\regs[30][12]~q ) # ((!dcifimemload_24)))) # (!\Mux19~2_combout  & (((\regs[26][12]~q  & dcifimemload_24))))

	.dataa(\regs[30][12]~q ),
	.datab(\regs[26][12]~q ),
	.datac(\Mux19~2_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hACF0;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N30
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\regs[20][12]~q ))) # (!dcifimemload_23 & (\regs[16][12]~q ))))

	.dataa(dcifimemload_24),
	.datab(\regs[16][12]~q ),
	.datac(\regs[20][12]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hFA44;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N14
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (dcifimemload_24 & ((\Mux19~4_combout  & ((\regs[28][12]~q ))) # (!\Mux19~4_combout  & (\regs[24][12]~q )))) # (!dcifimemload_24 & (((\Mux19~4_combout ))))

	.dataa(\regs[24][12]~q ),
	.datab(\regs[28][12]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux19~4_combout ),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hCFA0;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N8
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// \Mux19~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux19~3_combout )) # (!dcifimemload_22 & ((\Mux19~5_combout )))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux19~3_combout ),
	.datad(\Mux19~5_combout ),
	.cin(gnd),
	.combout(\Mux19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'hD9C8;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N4
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// \Mux19~7_combout  = (dcifimemload_24 & (((\regs[27][12]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[19][12]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[19][12]~q ),
	.datac(\regs[27][12]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hAAE4;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N26
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (dcifimemload_23 & ((\Mux19~7_combout  & (\regs[31][12]~q )) # (!\Mux19~7_combout  & ((\regs[23][12]~q ))))) # (!dcifimemload_23 & (((\Mux19~7_combout ))))

	.dataa(\regs[31][12]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[23][12]~q ),
	.datad(\Mux19~7_combout ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'hBBC0;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N14
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// \Mux19~9_combout  = (dcifimemload_21 & ((\Mux19~6_combout  & ((\Mux19~8_combout ))) # (!\Mux19~6_combout  & (\Mux19~1_combout )))) # (!dcifimemload_21 & (((\Mux19~6_combout ))))

	.dataa(\Mux19~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux19~6_combout ),
	.datad(\Mux19~8_combout ),
	.cin(gnd),
	.combout(\Mux19~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hF838;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N5
dffeas \regs[5][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][12] .is_wysiwyg = "true";
defparam \regs[5][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N4
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\regs[5][12]~q ))) # (!dcifimemload_21 & (\regs[4][12]~q ))))

	.dataa(dcifimemload_22),
	.datab(\regs[4][12]~q ),
	.datac(\regs[5][12]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hFA44;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N30
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (dcifimemload_22 & ((\Mux19~10_combout  & ((\regs[7][12]~q ))) # (!\Mux19~10_combout  & (\regs[6][12]~q )))) # (!dcifimemload_22 & (\Mux19~10_combout ))

	.dataa(dcifimemload_22),
	.datab(\Mux19~10_combout ),
	.datac(\regs[6][12]~q ),
	.datad(\regs[7][12]~q ),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hEC64;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N12
cycloneive_lcell_comb \Mux19~17 (
// Equation(s):
// \Mux19~17_combout  = (dcifimemload_21 & (((\regs[13][12]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][12]~q  & ((!dcifimemload_22))))

	.dataa(\regs[12][12]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[13][12]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux19~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~17 .lut_mask = 16'hCCE2;
defparam \Mux19~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N8
cycloneive_lcell_comb \Mux19~18 (
// Equation(s):
// \Mux19~18_combout  = (dcifimemload_22 & ((\Mux19~17_combout  & (\regs[15][12]~q )) # (!\Mux19~17_combout  & ((\regs[14][12]~q ))))) # (!dcifimemload_22 & (((\Mux19~17_combout ))))

	.dataa(\regs[15][12]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[14][12]~q ),
	.datad(\Mux19~17_combout ),
	.cin(gnd),
	.combout(\Mux19~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~18 .lut_mask = 16'hBBC0;
defparam \Mux19~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// \Mux19~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][12]~q ))) # (!dcifimemload_22 & (\regs[8][12]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][12]~q ),
	.datac(\regs[10][12]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux19~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hFA44;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N6
cycloneive_lcell_comb \Mux19~13 (
// Equation(s):
// \Mux19~13_combout  = (dcifimemload_21 & ((\Mux19~12_combout  & (\regs[11][12]~q )) # (!\Mux19~12_combout  & ((\regs[9][12]~q ))))) # (!dcifimemload_21 & (((\Mux19~12_combout ))))

	.dataa(\regs[11][12]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[9][12]~q ),
	.datad(\Mux19~12_combout ),
	.cin(gnd),
	.combout(\Mux19~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~13 .lut_mask = 16'hBBC0;
defparam \Mux19~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N29
dffeas \regs[3][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~38_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][12] .is_wysiwyg = "true";
defparam \regs[3][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N26
cycloneive_lcell_comb \Mux19~14 (
// Equation(s):
// \Mux19~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][12]~q ))) # (!dcifimemload_22 & (\regs[1][12]~q ))))

	.dataa(\regs[1][12]~q ),
	.datab(\regs[3][12]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux19~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~14 .lut_mask = 16'hC0A0;
defparam \Mux19~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N28
cycloneive_lcell_comb \Mux19~15 (
// Equation(s):
// \Mux19~15_combout  = (\Mux19~14_combout ) # ((\regs[2][12]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\regs[2][12]~q ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux19~14_combout ),
	.cin(gnd),
	.combout(\Mux19~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~15 .lut_mask = 16'hFF08;
defparam \Mux19~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N10
cycloneive_lcell_comb \Mux19~16 (
// Equation(s):
// \Mux19~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & (\Mux19~13_combout )) # (!dcifimemload_24 & ((\Mux19~15_combout )))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux19~13_combout ),
	.datad(\Mux19~15_combout ),
	.cin(gnd),
	.combout(\Mux19~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~16 .lut_mask = 16'hD9C8;
defparam \Mux19~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N24
cycloneive_lcell_comb \Mux19~19 (
// Equation(s):
// \Mux19~19_combout  = (dcifimemload_23 & ((\Mux19~16_combout  & ((\Mux19~18_combout ))) # (!\Mux19~16_combout  & (\Mux19~11_combout )))) # (!dcifimemload_23 & (((\Mux19~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux19~11_combout ),
	.datac(\Mux19~18_combout ),
	.datad(\Mux19~16_combout ),
	.cin(gnd),
	.combout(\Mux19~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~19 .lut_mask = 16'hF588;
defparam \Mux19~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N22
cycloneive_lcell_comb \regs~39 (
// Equation(s):
// \regs~39_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_11)) # (!cuifRegSel_0 & ((Mux203)))))

	.dataa(cuifRegSel_0),
	.datab(ramiframload_11),
	.datac(Mux201),
	.datad(cuifRegSel_11),
	.cin(gnd),
	.combout(\regs~39_combout ),
	.cout());
// synopsys translate_off
defparam \regs~39 .lut_mask = 16'h00D8;
defparam \regs~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N8
cycloneive_lcell_comb \regs~40 (
// Equation(s):
// \regs~40_combout  = (!\Equal0~1_combout  & ((\regs~39_combout ) # ((\Add1~18_combout  & \regs~64_combout ))))

	.dataa(\Equal0~1_combout ),
	.datab(Add19),
	.datac(\regs~39_combout ),
	.datad(\regs~64_combout ),
	.cin(gnd),
	.combout(\regs~40_combout ),
	.cout());
// synopsys translate_off
defparam \regs~40 .lut_mask = 16'h5450;
defparam \regs~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N20
cycloneive_lcell_comb \regs[23][11]~feeder (
// Equation(s):
// \regs[23][11]~feeder_combout  = \regs~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~40_combout ),
	.cin(gnd),
	.combout(\regs[23][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N21
dffeas \regs[23][11] (
	.clk(CLK),
	.d(\regs[23][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][11] .is_wysiwyg = "true";
defparam \regs[23][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N1
dffeas \regs[19][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][11] .is_wysiwyg = "true";
defparam \regs[19][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N13
dffeas \regs[27][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][11] .is_wysiwyg = "true";
defparam \regs[27][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N12
cycloneive_lcell_comb \Mux52~7 (
// Equation(s):
// \Mux52~7_combout  = (dcifimemload_19 & (((\regs[27][11]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\regs[19][11]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\regs[19][11]~q ),
	.datac(\regs[27][11]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux52~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~7 .lut_mask = 16'hAAE4;
defparam \Mux52~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N15
dffeas \regs[31][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][11] .is_wysiwyg = "true";
defparam \regs[31][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N10
cycloneive_lcell_comb \Mux52~8 (
// Equation(s):
// \Mux52~8_combout  = (dcifimemload_18 & ((\Mux52~7_combout  & ((\regs[31][11]~q ))) # (!\Mux52~7_combout  & (\regs[23][11]~q )))) # (!dcifimemload_18 & (((\Mux52~7_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[23][11]~q ),
	.datac(\Mux52~7_combout ),
	.datad(\regs[31][11]~q ),
	.cin(gnd),
	.combout(\Mux52~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~8 .lut_mask = 16'hF858;
defparam \Mux52~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N9
dffeas \regs[29][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][11] .is_wysiwyg = "true";
defparam \regs[29][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N28
cycloneive_lcell_comb \regs[21][11]~feeder (
// Equation(s):
// \regs[21][11]~feeder_combout  = \regs~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~40_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[21][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][11]~feeder .lut_mask = 16'hF0F0;
defparam \regs[21][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N29
dffeas \regs[21][11] (
	.clk(CLK),
	.d(\regs[21][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][11] .is_wysiwyg = "true";
defparam \regs[21][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N30
cycloneive_lcell_comb \regs[25][11]~feeder (
// Equation(s):
// \regs[25][11]~feeder_combout  = \regs~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~40_combout ),
	.cin(gnd),
	.combout(\regs[25][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[25][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[25][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N31
dffeas \regs[25][11] (
	.clk(CLK),
	.d(\regs[25][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][11] .is_wysiwyg = "true";
defparam \regs[25][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N2
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (dcifimemload_19 & (((\regs[25][11]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\regs[17][11]~q  & ((!dcifimemload_18))))

	.dataa(\regs[17][11]~q ),
	.datab(\regs[25][11]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hF0CA;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N8
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (dcifimemload_18 & ((\Mux52~0_combout  & (\regs[29][11]~q )) # (!\Mux52~0_combout  & ((\regs[21][11]~q ))))) # (!dcifimemload_18 & (((\Mux52~0_combout ))))

	.dataa(\regs[29][11]~q ),
	.datab(\regs[21][11]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux52~0_combout ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hAFC0;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N17
dffeas \regs[20][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][11] .is_wysiwyg = "true";
defparam \regs[20][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N16
cycloneive_lcell_comb \Mux52~4 (
// Equation(s):
// \Mux52~4_combout  = (dcifimemload_18 & (((\regs[20][11]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[16][11]~q  & ((!dcifimemload_19))))

	.dataa(\regs[16][11]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[20][11]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux52~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~4 .lut_mask = 16'hCCE2;
defparam \Mux52~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N15
dffeas \regs[24][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][11] .is_wysiwyg = "true";
defparam \regs[24][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N14
cycloneive_lcell_comb \Mux52~5 (
// Equation(s):
// \Mux52~5_combout  = (\Mux52~4_combout  & ((\regs[28][11]~q ) # ((!dcifimemload_19)))) # (!\Mux52~4_combout  & (((\regs[24][11]~q  & dcifimemload_19))))

	.dataa(\regs[28][11]~q ),
	.datab(\Mux52~4_combout ),
	.datac(\regs[24][11]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux52~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~5 .lut_mask = 16'hB8CC;
defparam \Mux52~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N14
cycloneive_lcell_comb \regs[26][11]~feeder (
// Equation(s):
// \regs[26][11]~feeder_combout  = \regs~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~40_combout ),
	.cin(gnd),
	.combout(\regs[26][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[26][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N15
dffeas \regs[26][11] (
	.clk(CLK),
	.d(\regs[26][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][11] .is_wysiwyg = "true";
defparam \regs[26][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N9
dffeas \regs[22][11] (
	.clk(CLK),
	.d(\regs~40_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][11] .is_wysiwyg = "true";
defparam \regs[22][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N8
cycloneive_lcell_comb \Mux52~2 (
// Equation(s):
// \Mux52~2_combout  = (dcifimemload_18 & (((\regs[22][11]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[18][11]~q  & ((!dcifimemload_19))))

	.dataa(\regs[18][11]~q ),
	.datab(\regs[22][11]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux52~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~2 .lut_mask = 16'hF0CA;
defparam \Mux52~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N28
cycloneive_lcell_comb \Mux52~3 (
// Equation(s):
// \Mux52~3_combout  = (\Mux52~2_combout  & ((\regs[30][11]~q ) # ((!dcifimemload_19)))) # (!\Mux52~2_combout  & (((\regs[26][11]~q  & dcifimemload_19))))

	.dataa(\regs[30][11]~q ),
	.datab(\regs[26][11]~q ),
	.datac(\Mux52~2_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux52~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~3 .lut_mask = 16'hACF0;
defparam \Mux52~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N2
cycloneive_lcell_comb \Mux52~6 (
// Equation(s):
// \Mux52~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux52~3_combout ))) # (!dcifimemload_17 & (\Mux52~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux52~5_combout ),
	.datad(\Mux52~3_combout ),
	.cin(gnd),
	.combout(\Mux52~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~6 .lut_mask = 16'hDC98;
defparam \Mux52~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N13
dffeas \regs[14][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][11] .is_wysiwyg = "true";
defparam \regs[14][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N4
cycloneive_lcell_comb \regs[15][11]~feeder (
// Equation(s):
// \regs[15][11]~feeder_combout  = \regs~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~40_combout ),
	.cin(gnd),
	.combout(\regs[15][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N5
dffeas \regs[15][11] (
	.clk(CLK),
	.d(\regs[15][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][11] .is_wysiwyg = "true";
defparam \regs[15][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y44_N5
dffeas \regs[12][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][11] .is_wysiwyg = "true";
defparam \regs[12][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N4
cycloneive_lcell_comb \Mux52~17 (
// Equation(s):
// \Mux52~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][11]~q )) # (!dcifimemload_16 & ((\regs[12][11]~q )))))

	.dataa(\regs[13][11]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][11]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux52~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~17 .lut_mask = 16'hEE30;
defparam \Mux52~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N14
cycloneive_lcell_comb \Mux52~18 (
// Equation(s):
// \Mux52~18_combout  = (\Mux52~17_combout  & (((\regs[15][11]~q ) # (!dcifimemload_17)))) # (!\Mux52~17_combout  & (\regs[14][11]~q  & ((dcifimemload_17))))

	.dataa(\regs[14][11]~q ),
	.datab(\regs[15][11]~q ),
	.datac(\Mux52~17_combout ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux52~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~18 .lut_mask = 16'hCAF0;
defparam \Mux52~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N31
dffeas \regs[2][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][11] .is_wysiwyg = "true";
defparam \regs[2][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N15
dffeas \regs[3][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][11] .is_wysiwyg = "true";
defparam \regs[3][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N13
dffeas \regs[1][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][11] .is_wysiwyg = "true";
defparam \regs[1][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N12
cycloneive_lcell_comb \Mux52~14 (
// Equation(s):
// \Mux52~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][11]~q )) # (!dcifimemload_17 & ((\regs[1][11]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[3][11]~q ),
	.datac(\regs[1][11]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux52~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~14 .lut_mask = 16'hD800;
defparam \Mux52~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N30
cycloneive_lcell_comb \Mux52~15 (
// Equation(s):
// \Mux52~15_combout  = (\Mux52~14_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][11]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[2][11]~q ),
	.datad(\Mux52~14_combout ),
	.cin(gnd),
	.combout(\Mux52~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~15 .lut_mask = 16'hFF20;
defparam \Mux52~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N22
cycloneive_lcell_comb \regs[9][11]~feeder (
// Equation(s):
// \regs[9][11]~feeder_combout  = \regs~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~40_combout ),
	.cin(gnd),
	.combout(\regs[9][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N23
dffeas \regs[9][11] (
	.clk(CLK),
	.d(\regs[9][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][11] .is_wysiwyg = "true";
defparam \regs[9][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N7
dffeas \regs[11][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][11] .is_wysiwyg = "true";
defparam \regs[11][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N21
dffeas \regs[10][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][11] .is_wysiwyg = "true";
defparam \regs[10][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N17
dffeas \regs[8][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][11] .is_wysiwyg = "true";
defparam \regs[8][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N16
cycloneive_lcell_comb \Mux52~12 (
// Equation(s):
// \Mux52~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][11]~q )) # (!dcifimemload_17 & ((\regs[8][11]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][11]~q ),
	.datac(\regs[8][11]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux52~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~12 .lut_mask = 16'hEE50;
defparam \Mux52~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N6
cycloneive_lcell_comb \Mux52~13 (
// Equation(s):
// \Mux52~13_combout  = (dcifimemload_16 & ((\Mux52~12_combout  & ((\regs[11][11]~q ))) # (!\Mux52~12_combout  & (\regs[9][11]~q )))) # (!dcifimemload_16 & (((\Mux52~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][11]~q ),
	.datac(\regs[11][11]~q ),
	.datad(\Mux52~12_combout ),
	.cin(gnd),
	.combout(\Mux52~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~13 .lut_mask = 16'hF588;
defparam \Mux52~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N26
cycloneive_lcell_comb \Mux52~16 (
// Equation(s):
// \Mux52~16_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux52~13_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & (\Mux52~15_combout )))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux52~15_combout ),
	.datad(\Mux52~13_combout ),
	.cin(gnd),
	.combout(\Mux52~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~16 .lut_mask = 16'hBA98;
defparam \Mux52~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N7
dffeas \regs[7][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][11] .is_wysiwyg = "true";
defparam \regs[7][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N15
dffeas \regs[5][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][11] .is_wysiwyg = "true";
defparam \regs[5][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N14
cycloneive_lcell_comb \Mux52~10 (
// Equation(s):
// \Mux52~10_combout  = (dcifimemload_16 & (((\regs[5][11]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][11]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][11]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[5][11]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux52~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~10 .lut_mask = 16'hCCE2;
defparam \Mux52~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N21
dffeas \regs[6][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][11] .is_wysiwyg = "true";
defparam \regs[6][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N20
cycloneive_lcell_comb \Mux52~11 (
// Equation(s):
// \Mux52~11_combout  = (\Mux52~10_combout  & ((\regs[7][11]~q ) # ((!dcifimemload_17)))) # (!\Mux52~10_combout  & (((\regs[6][11]~q  & dcifimemload_17))))

	.dataa(\regs[7][11]~q ),
	.datab(\Mux52~10_combout ),
	.datac(\regs[6][11]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux52~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~11 .lut_mask = 16'hB8CC;
defparam \Mux52~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N17
dffeas \regs[4][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][11] .is_wysiwyg = "true";
defparam \regs[4][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N16
cycloneive_lcell_comb \Mux20~12 (
// Equation(s):
// \Mux20~12_combout  = (dcifimemload_21 & ((\regs[5][11]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\regs[4][11]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[5][11]~q ),
	.datac(\regs[4][11]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux20~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~12 .lut_mask = 16'hAAD8;
defparam \Mux20~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N6
cycloneive_lcell_comb \Mux20~13 (
// Equation(s):
// \Mux20~13_combout  = (dcifimemload_22 & ((\Mux20~12_combout  & ((\regs[7][11]~q ))) # (!\Mux20~12_combout  & (\regs[6][11]~q )))) # (!dcifimemload_22 & (((\Mux20~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[6][11]~q ),
	.datac(\regs[7][11]~q ),
	.datad(\Mux20~12_combout ),
	.cin(gnd),
	.combout(\Mux20~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~13 .lut_mask = 16'hF588;
defparam \Mux20~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N14
cycloneive_lcell_comb \Mux20~14 (
// Equation(s):
// \Mux20~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][11]~q ))) # (!dcifimemload_22 & (\regs[1][11]~q ))))

	.dataa(\regs[1][11]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[3][11]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux20~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~14 .lut_mask = 16'hC088;
defparam \Mux20~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N24
cycloneive_lcell_comb \Mux20~15 (
// Equation(s):
// \Mux20~15_combout  = (\Mux20~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][11]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[2][11]~q ),
	.datad(\Mux20~14_combout ),
	.cin(gnd),
	.combout(\Mux20~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~15 .lut_mask = 16'hFF20;
defparam \Mux20~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N26
cycloneive_lcell_comb \Mux20~16 (
// Equation(s):
// \Mux20~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux20~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & ((\Mux20~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux20~13_combout ),
	.datad(\Mux20~15_combout ),
	.cin(gnd),
	.combout(\Mux20~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~16 .lut_mask = 16'hB9A8;
defparam \Mux20~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N12
cycloneive_lcell_comb \Mux20~18 (
// Equation(s):
// \Mux20~18_combout  = (\Mux20~17_combout  & ((\regs[15][11]~q ) # ((!dcifimemload_22)))) # (!\Mux20~17_combout  & (((\regs[14][11]~q  & dcifimemload_22))))

	.dataa(\Mux20~17_combout ),
	.datab(\regs[15][11]~q ),
	.datac(\regs[14][11]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux20~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~18 .lut_mask = 16'hD8AA;
defparam \Mux20~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N20
cycloneive_lcell_comb \Mux20~10 (
// Equation(s):
// \Mux20~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][11]~q ))) # (!dcifimemload_22 & (\regs[8][11]~q ))))

	.dataa(\regs[8][11]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[10][11]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux20~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~10 .lut_mask = 16'hFC22;
defparam \Mux20~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N24
cycloneive_lcell_comb \Mux20~11 (
// Equation(s):
// \Mux20~11_combout  = (\Mux20~10_combout  & (((\regs[11][11]~q ) # (!dcifimemload_21)))) # (!\Mux20~10_combout  & (\regs[9][11]~q  & ((dcifimemload_21))))

	.dataa(\regs[9][11]~q ),
	.datab(\regs[11][11]~q ),
	.datac(\Mux20~10_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux20~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~11 .lut_mask = 16'hCAF0;
defparam \Mux20~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N8
cycloneive_lcell_comb \Mux20~19 (
// Equation(s):
// \Mux20~19_combout  = (\Mux20~16_combout  & (((\Mux20~18_combout )) # (!dcifimemload_24))) # (!\Mux20~16_combout  & (dcifimemload_24 & ((\Mux20~11_combout ))))

	.dataa(\Mux20~16_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux20~18_combout ),
	.datad(\Mux20~11_combout ),
	.cin(gnd),
	.combout(\Mux20~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~19 .lut_mask = 16'hE6A2;
defparam \Mux20~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N0
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// \Mux20~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[23][11]~q )) # (!dcifimemload_23 & ((\regs[19][11]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[23][11]~q ),
	.datac(\regs[19][11]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hEE50;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N14
cycloneive_lcell_comb \Mux20~8 (
// Equation(s):
// \Mux20~8_combout  = (dcifimemload_24 & ((\Mux20~7_combout  & ((\regs[31][11]~q ))) # (!\Mux20~7_combout  & (\regs[27][11]~q )))) # (!dcifimemload_24 & (((\Mux20~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][11]~q ),
	.datac(\regs[31][11]~q ),
	.datad(\Mux20~7_combout ),
	.cin(gnd),
	.combout(\Mux20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~8 .lut_mask = 16'hF588;
defparam \Mux20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N30
cycloneive_lcell_comb \regs[17][11]~feeder (
// Equation(s):
// \regs[17][11]~feeder_combout  = \regs~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~40_combout ),
	.cin(gnd),
	.combout(\regs[17][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[17][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N31
dffeas \regs[17][11] (
	.clk(CLK),
	.d(\regs[17][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][11] .is_wysiwyg = "true";
defparam \regs[17][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N14
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[21][11]~q )) # (!dcifimemload_23 & ((\regs[17][11]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[21][11]~q ),
	.datac(\regs[17][11]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hEE50;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N8
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (dcifimemload_24 & ((\Mux20~0_combout  & (\regs[29][11]~q )) # (!\Mux20~0_combout  & ((\regs[25][11]~q ))))) # (!dcifimemload_24 & (\Mux20~0_combout ))

	.dataa(dcifimemload_24),
	.datab(\Mux20~0_combout ),
	.datac(\regs[29][11]~q ),
	.datad(\regs[25][11]~q ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hE6C4;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N7
dffeas \regs[28][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][11] .is_wysiwyg = "true";
defparam \regs[28][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N17
dffeas \regs[16][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~40_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][11] .is_wysiwyg = "true";
defparam \regs[16][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N16
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[24][11]~q )) # (!dcifimemload_24 & ((\regs[16][11]~q )))))

	.dataa(dcifimemload_23),
	.datab(\regs[24][11]~q ),
	.datac(\regs[16][11]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hEE50;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N6
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// \Mux20~5_combout  = (dcifimemload_23 & ((\Mux20~4_combout  & ((\regs[28][11]~q ))) # (!\Mux20~4_combout  & (\regs[20][11]~q )))) # (!dcifimemload_23 & (((\Mux20~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[20][11]~q ),
	.datac(\regs[28][11]~q ),
	.datad(\Mux20~4_combout ),
	.cin(gnd),
	.combout(\Mux20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hF588;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N8
cycloneive_lcell_comb \regs[18][11]~feeder (
// Equation(s):
// \regs[18][11]~feeder_combout  = \regs~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~40_combout ),
	.cin(gnd),
	.combout(\regs[18][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[18][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[18][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N9
dffeas \regs[18][11] (
	.clk(CLK),
	.d(\regs[18][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][11] .is_wysiwyg = "true";
defparam \regs[18][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N16
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (dcifimemload_24 & ((\regs[26][11]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[18][11]~q  & !dcifimemload_23))))

	.dataa(\regs[26][11]~q ),
	.datab(\regs[18][11]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hF0AC;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N14
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (dcifimemload_23 & ((\Mux20~2_combout  & (\regs[30][11]~q )) # (!\Mux20~2_combout  & ((\regs[22][11]~q ))))) # (!dcifimemload_23 & (((\Mux20~2_combout ))))

	.dataa(\regs[30][11]~q ),
	.datab(\regs[22][11]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux20~2_combout ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hAFC0;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N20
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// \Mux20~6_combout  = (dcifimemload_22 & (((dcifimemload_21) # (\Mux20~3_combout )))) # (!dcifimemload_22 & (\Mux20~5_combout  & (!dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\Mux20~5_combout ),
	.datac(dcifimemload_21),
	.datad(\Mux20~3_combout ),
	.cin(gnd),
	.combout(\Mux20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'hAEA4;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N2
cycloneive_lcell_comb \Mux20~9 (
// Equation(s):
// \Mux20~9_combout  = (dcifimemload_21 & ((\Mux20~6_combout  & (\Mux20~8_combout )) # (!\Mux20~6_combout  & ((\Mux20~1_combout ))))) # (!dcifimemload_21 & (((\Mux20~6_combout ))))

	.dataa(\Mux20~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux20~1_combout ),
	.datad(\Mux20~6_combout ),
	.cin(gnd),
	.combout(\Mux20~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~9 .lut_mask = 16'hBBC0;
defparam \Mux20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N0
cycloneive_lcell_comb \regs~41 (
// Equation(s):
// \regs~41_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_10)) # (!cuifRegSel_0 & ((Mux213)))))

	.dataa(cuifRegSel_0),
	.datab(cuifRegSel_11),
	.datac(ramiframload_10),
	.datad(Mux211),
	.cin(gnd),
	.combout(\regs~41_combout ),
	.cout());
// synopsys translate_off
defparam \regs~41 .lut_mask = 16'h3120;
defparam \regs~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N14
cycloneive_lcell_comb \regs~42 (
// Equation(s):
// \regs~42_combout  = (!\Equal0~1_combout  & ((\regs~41_combout ) # ((\regs~64_combout  & \Add1~16_combout ))))

	.dataa(\regs~64_combout ),
	.datab(Add18),
	.datac(\Equal0~1_combout ),
	.datad(\regs~41_combout ),
	.cin(gnd),
	.combout(\regs~42_combout ),
	.cout());
// synopsys translate_off
defparam \regs~42 .lut_mask = 16'h0F08;
defparam \regs~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N1
dffeas \regs[27][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][10] .is_wysiwyg = "true";
defparam \regs[27][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N7
dffeas \regs[31][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][10] .is_wysiwyg = "true";
defparam \regs[31][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N4
cycloneive_lcell_comb \regs[19][10]~feeder (
// Equation(s):
// \regs[19][10]~feeder_combout  = \regs~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~42_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[19][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][10]~feeder .lut_mask = 16'hF0F0;
defparam \regs[19][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N5
dffeas \regs[19][10] (
	.clk(CLK),
	.d(\regs[19][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][10] .is_wysiwyg = "true";
defparam \regs[19][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N4
cycloneive_lcell_comb \Mux53~7 (
// Equation(s):
// \Mux53~7_combout  = (dcifimemload_18 & ((\regs[23][10]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[19][10]~q  & !dcifimemload_19))))

	.dataa(\regs[23][10]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[19][10]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux53~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~7 .lut_mask = 16'hCCB8;
defparam \Mux53~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N22
cycloneive_lcell_comb \Mux53~8 (
// Equation(s):
// \Mux53~8_combout  = (\Mux53~7_combout  & (((\regs[31][10]~q ) # (!dcifimemload_19)))) # (!\Mux53~7_combout  & (\regs[27][10]~q  & ((dcifimemload_19))))

	.dataa(\regs[27][10]~q ),
	.datab(\regs[31][10]~q ),
	.datac(\Mux53~7_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux53~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~8 .lut_mask = 16'hCAF0;
defparam \Mux53~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N31
dffeas \regs[30][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][10] .is_wysiwyg = "true";
defparam \regs[30][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N21
dffeas \regs[18][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][10] .is_wysiwyg = "true";
defparam \regs[18][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N16
cycloneive_lcell_comb \Mux53~2 (
// Equation(s):
// \Mux53~2_combout  = (dcifimemload_19 & ((\regs[26][10]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\regs[18][10]~q  & !dcifimemload_18))))

	.dataa(\regs[26][10]~q ),
	.datab(\regs[18][10]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux53~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~2 .lut_mask = 16'hF0AC;
defparam \Mux53~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N6
cycloneive_lcell_comb \Mux53~3 (
// Equation(s):
// \Mux53~3_combout  = (dcifimemload_18 & ((\Mux53~2_combout  & ((\regs[30][10]~q ))) # (!\Mux53~2_combout  & (\regs[22][10]~q )))) # (!dcifimemload_18 & (((\Mux53~2_combout ))))

	.dataa(\regs[22][10]~q ),
	.datab(\regs[30][10]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux53~2_combout ),
	.cin(gnd),
	.combout(\Mux53~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~3 .lut_mask = 16'hCFA0;
defparam \Mux53~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N23
dffeas \regs[28][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][10] .is_wysiwyg = "true";
defparam \regs[28][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N7
dffeas \regs[20][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][10] .is_wysiwyg = "true";
defparam \regs[20][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N3
dffeas \regs[24][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][10] .is_wysiwyg = "true";
defparam \regs[24][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N2
cycloneive_lcell_comb \Mux53~4 (
// Equation(s):
// \Mux53~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[24][10]~q ))) # (!dcifimemload_19 & (\regs[16][10]~q ))))

	.dataa(\regs[16][10]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[24][10]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux53~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~4 .lut_mask = 16'hFC22;
defparam \Mux53~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N6
cycloneive_lcell_comb \Mux53~5 (
// Equation(s):
// \Mux53~5_combout  = (dcifimemload_18 & ((\Mux53~4_combout  & (\regs[28][10]~q )) # (!\Mux53~4_combout  & ((\regs[20][10]~q ))))) # (!dcifimemload_18 & (((\Mux53~4_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[28][10]~q ),
	.datac(\regs[20][10]~q ),
	.datad(\Mux53~4_combout ),
	.cin(gnd),
	.combout(\Mux53~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~5 .lut_mask = 16'hDDA0;
defparam \Mux53~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N4
cycloneive_lcell_comb \Mux53~6 (
// Equation(s):
// \Mux53~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux53~3_combout )) # (!dcifimemload_17 & ((\Mux53~5_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux53~3_combout ),
	.datad(\Mux53~5_combout ),
	.cin(gnd),
	.combout(\Mux53~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~6 .lut_mask = 16'hD9C8;
defparam \Mux53~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N28
cycloneive_lcell_comb \regs[29][10]~feeder (
// Equation(s):
// \regs[29][10]~feeder_combout  = \regs~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~42_combout ),
	.cin(gnd),
	.combout(\regs[29][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][10]~feeder .lut_mask = 16'hFF00;
defparam \regs[29][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y45_N29
dffeas \regs[29][10] (
	.clk(CLK),
	.d(\regs[29][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][10] .is_wysiwyg = "true";
defparam \regs[29][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N3
dffeas \regs[25][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][10] .is_wysiwyg = "true";
defparam \regs[25][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N31
dffeas \regs[21][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][10] .is_wysiwyg = "true";
defparam \regs[21][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N30
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (dcifimemload_18 & (((\regs[21][10]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[17][10]~q  & ((!dcifimemload_19))))

	.dataa(\regs[17][10]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[21][10]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hCCE2;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N2
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (dcifimemload_19 & ((\Mux53~0_combout  & (\regs[29][10]~q )) # (!\Mux53~0_combout  & ((\regs[25][10]~q ))))) # (!dcifimemload_19 & (((\Mux53~0_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[29][10]~q ),
	.datac(\regs[25][10]~q ),
	.datad(\Mux53~0_combout ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hDDA0;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N13
dffeas \regs[14][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][10] .is_wysiwyg = "true";
defparam \regs[14][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N3
dffeas \regs[15][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][10] .is_wysiwyg = "true";
defparam \regs[15][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N5
dffeas \regs[13][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][10] .is_wysiwyg = "true";
defparam \regs[13][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N31
dffeas \regs[12][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][10] .is_wysiwyg = "true";
defparam \regs[12][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N30
cycloneive_lcell_comb \Mux53~17 (
// Equation(s):
// \Mux53~17_combout  = (dcifimemload_16 & ((\regs[13][10]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[12][10]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[13][10]~q ),
	.datac(\regs[12][10]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux53~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~17 .lut_mask = 16'hAAD8;
defparam \Mux53~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N2
cycloneive_lcell_comb \Mux53~18 (
// Equation(s):
// \Mux53~18_combout  = (dcifimemload_17 & ((\Mux53~17_combout  & ((\regs[15][10]~q ))) # (!\Mux53~17_combout  & (\regs[14][10]~q )))) # (!dcifimemload_17 & (((\Mux53~17_combout ))))

	.dataa(\regs[14][10]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[15][10]~q ),
	.datad(\Mux53~17_combout ),
	.cin(gnd),
	.combout(\Mux53~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~18 .lut_mask = 16'hF388;
defparam \Mux53~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N13
dffeas \regs[11][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][10] .is_wysiwyg = "true";
defparam \regs[11][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N15
dffeas \regs[10][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][10] .is_wysiwyg = "true";
defparam \regs[10][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N14
cycloneive_lcell_comb \Mux53~10 (
// Equation(s):
// \Mux53~10_combout  = (dcifimemload_17 & (((\regs[10][10]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\regs[8][10]~q  & ((!dcifimemload_16))))

	.dataa(\regs[8][10]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[10][10]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux53~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~10 .lut_mask = 16'hCCE2;
defparam \Mux53~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N13
dffeas \regs[9][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][10] .is_wysiwyg = "true";
defparam \regs[9][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N12
cycloneive_lcell_comb \Mux53~11 (
// Equation(s):
// \Mux53~11_combout  = (\Mux53~10_combout  & ((\regs[11][10]~q ) # ((!dcifimemload_16)))) # (!\Mux53~10_combout  & (((\regs[9][10]~q  & dcifimemload_16))))

	.dataa(\regs[11][10]~q ),
	.datab(\Mux53~10_combout ),
	.datac(\regs[9][10]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux53~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~11 .lut_mask = 16'hB8CC;
defparam \Mux53~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y45_N7
dffeas \regs[2][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][10] .is_wysiwyg = "true";
defparam \regs[2][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y45_N21
dffeas \regs[1][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][10] .is_wysiwyg = "true";
defparam \regs[1][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N20
cycloneive_lcell_comb \Mux53~14 (
// Equation(s):
// \Mux53~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][10]~q )) # (!dcifimemload_17 & ((\regs[1][10]~q )))))

	.dataa(\regs[3][10]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[1][10]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux53~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~14 .lut_mask = 16'hB800;
defparam \Mux53~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N6
cycloneive_lcell_comb \Mux53~15 (
// Equation(s):
// \Mux53~15_combout  = (\Mux53~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][10]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][10]~q ),
	.datad(\Mux53~14_combout ),
	.cin(gnd),
	.combout(\Mux53~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~15 .lut_mask = 16'hFF40;
defparam \Mux53~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N17
dffeas \regs[7][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][10] .is_wysiwyg = "true";
defparam \regs[7][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N14
cycloneive_lcell_comb \regs[5][10]~feeder (
// Equation(s):
// \regs[5][10]~feeder_combout  = \regs~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~42_combout ),
	.cin(gnd),
	.combout(\regs[5][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][10]~feeder .lut_mask = 16'hFF00;
defparam \regs[5][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y45_N15
dffeas \regs[5][10] (
	.clk(CLK),
	.d(\regs[5][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][10] .is_wysiwyg = "true";
defparam \regs[5][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N5
dffeas \regs[4][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][10] .is_wysiwyg = "true";
defparam \regs[4][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N4
cycloneive_lcell_comb \Mux53~12 (
// Equation(s):
// \Mux53~12_combout  = (dcifimemload_16 & ((\regs[5][10]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][10]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[5][10]~q ),
	.datac(\regs[4][10]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux53~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~12 .lut_mask = 16'hAAD8;
defparam \Mux53~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N16
cycloneive_lcell_comb \Mux53~13 (
// Equation(s):
// \Mux53~13_combout  = (dcifimemload_17 & ((\Mux53~12_combout  & ((\regs[7][10]~q ))) # (!\Mux53~12_combout  & (\regs[6][10]~q )))) # (!dcifimemload_17 & (((\Mux53~12_combout ))))

	.dataa(\regs[6][10]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[7][10]~q ),
	.datad(\Mux53~12_combout ),
	.cin(gnd),
	.combout(\Mux53~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~13 .lut_mask = 16'hF388;
defparam \Mux53~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N0
cycloneive_lcell_comb \Mux53~16 (
// Equation(s):
// \Mux53~16_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux53~13_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & (\Mux53~15_combout )))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux53~15_combout ),
	.datad(\Mux53~13_combout ),
	.cin(gnd),
	.combout(\Mux53~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~16 .lut_mask = 16'hBA98;
defparam \Mux53~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N3
dffeas \regs[23][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][10] .is_wysiwyg = "true";
defparam \regs[23][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N0
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// \Mux21~7_combout  = (dcifimemload_24 & (((\regs[27][10]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[19][10]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[19][10]~q ),
	.datac(\regs[27][10]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hAAE4;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N6
cycloneive_lcell_comb \Mux21~8 (
// Equation(s):
// \Mux21~8_combout  = (dcifimemload_23 & ((\Mux21~7_combout  & ((\regs[31][10]~q ))) # (!\Mux21~7_combout  & (\regs[23][10]~q )))) # (!dcifimemload_23 & (((\Mux21~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[23][10]~q ),
	.datac(\regs[31][10]~q ),
	.datad(\Mux21~7_combout ),
	.cin(gnd),
	.combout(\Mux21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~8 .lut_mask = 16'hF588;
defparam \Mux21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N24
cycloneive_lcell_comb \regs[16][10]~feeder (
// Equation(s):
// \regs[16][10]~feeder_combout  = \regs~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~42_combout ),
	.cin(gnd),
	.combout(\regs[16][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[16][10]~feeder .lut_mask = 16'hFF00;
defparam \regs[16][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N25
dffeas \regs[16][10] (
	.clk(CLK),
	.d(\regs[16][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][10] .is_wysiwyg = "true";
defparam \regs[16][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N20
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (dcifimemload_23 & ((\regs[20][10]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[16][10]~q  & !dcifimemload_24))))

	.dataa(\regs[20][10]~q ),
	.datab(\regs[16][10]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hF0AC;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N22
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// \Mux21~5_combout  = (dcifimemload_24 & ((\Mux21~4_combout  & ((\regs[28][10]~q ))) # (!\Mux21~4_combout  & (\regs[24][10]~q )))) # (!dcifimemload_24 & (((\Mux21~4_combout ))))

	.dataa(\regs[24][10]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[28][10]~q ),
	.datad(\Mux21~4_combout ),
	.cin(gnd),
	.combout(\Mux21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hF388;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N4
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// \Mux21~6_combout  = (dcifimemload_22 & ((\Mux21~3_combout ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((!dcifimemload_21 & \Mux21~5_combout ))))

	.dataa(\Mux21~3_combout ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux21~5_combout ),
	.cin(gnd),
	.combout(\Mux21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'hCBC8;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N5
dffeas \regs[17][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][10] .is_wysiwyg = "true";
defparam \regs[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N4
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (dcifimemload_24 & ((\regs[25][10]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[17][10]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[25][10]~q ),
	.datac(\regs[17][10]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hAAD8;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N6
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (dcifimemload_23 & ((\Mux21~0_combout  & (\regs[29][10]~q )) # (!\Mux21~0_combout  & ((\regs[21][10]~q ))))) # (!dcifimemload_23 & (((\Mux21~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[29][10]~q ),
	.datac(\regs[21][10]~q ),
	.datad(\Mux21~0_combout ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hDDA0;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N30
cycloneive_lcell_comb \Mux21~9 (
// Equation(s):
// \Mux21~9_combout  = (dcifimemload_21 & ((\Mux21~6_combout  & (\Mux21~8_combout )) # (!\Mux21~6_combout  & ((\Mux21~1_combout ))))) # (!dcifimemload_21 & (((\Mux21~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux21~8_combout ),
	.datac(\Mux21~6_combout ),
	.datad(\Mux21~1_combout ),
	.cin(gnd),
	.combout(\Mux21~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~9 .lut_mask = 16'hDAD0;
defparam \Mux21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N12
cycloneive_lcell_comb \regs[6][10]~feeder (
// Equation(s):
// \regs[6][10]~feeder_combout  = \regs~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~42_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[6][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][10]~feeder .lut_mask = 16'hF0F0;
defparam \regs[6][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N13
dffeas \regs[6][10] (
	.clk(CLK),
	.d(\regs[6][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][10] .is_wysiwyg = "true";
defparam \regs[6][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N20
cycloneive_lcell_comb \Mux21~10 (
// Equation(s):
// \Mux21~10_combout  = (dcifimemload_21 & (((\regs[5][10]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][10]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][10]~q ),
	.datac(\regs[5][10]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux21~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~10 .lut_mask = 16'hAAE4;
defparam \Mux21~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y45_N22
cycloneive_lcell_comb \Mux21~11 (
// Equation(s):
// \Mux21~11_combout  = (dcifimemload_22 & ((\Mux21~10_combout  & (\regs[7][10]~q )) # (!\Mux21~10_combout  & ((\regs[6][10]~q ))))) # (!dcifimemload_22 & (((\Mux21~10_combout ))))

	.dataa(\regs[7][10]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[6][10]~q ),
	.datad(\Mux21~10_combout ),
	.cin(gnd),
	.combout(\Mux21~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~11 .lut_mask = 16'hBBC0;
defparam \Mux21~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N4
cycloneive_lcell_comb \Mux21~17 (
// Equation(s):
// \Mux21~17_combout  = (dcifimemload_21 & (((\regs[13][10]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][10]~q  & ((!dcifimemload_22))))

	.dataa(\regs[12][10]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[13][10]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux21~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~17 .lut_mask = 16'hCCE2;
defparam \Mux21~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N12
cycloneive_lcell_comb \Mux21~18 (
// Equation(s):
// \Mux21~18_combout  = (dcifimemload_22 & ((\Mux21~17_combout  & ((\regs[15][10]~q ))) # (!\Mux21~17_combout  & (\regs[14][10]~q )))) # (!dcifimemload_22 & (\Mux21~17_combout ))

	.dataa(dcifimemload_22),
	.datab(\Mux21~17_combout ),
	.datac(\regs[14][10]~q ),
	.datad(\regs[15][10]~q ),
	.cin(gnd),
	.combout(\Mux21~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~18 .lut_mask = 16'hEC64;
defparam \Mux21~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N3
dffeas \regs[8][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~42_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][10] .is_wysiwyg = "true";
defparam \regs[8][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N2
cycloneive_lcell_comb \Mux21~12 (
// Equation(s):
// \Mux21~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\regs[10][10]~q )) # (!dcifimemload_22 & ((\regs[8][10]~q )))))

	.dataa(\regs[10][10]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[8][10]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux21~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~12 .lut_mask = 16'hEE30;
defparam \Mux21~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N12
cycloneive_lcell_comb \Mux21~13 (
// Equation(s):
// \Mux21~13_combout  = (dcifimemload_21 & ((\Mux21~12_combout  & ((\regs[11][10]~q ))) # (!\Mux21~12_combout  & (\regs[9][10]~q )))) # (!dcifimemload_21 & (((\Mux21~12_combout ))))

	.dataa(\regs[9][10]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[11][10]~q ),
	.datad(\Mux21~12_combout ),
	.cin(gnd),
	.combout(\Mux21~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~13 .lut_mask = 16'hF388;
defparam \Mux21~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N10
cycloneive_lcell_comb \regs[3][10]~feeder (
// Equation(s):
// \regs[3][10]~feeder_combout  = \regs~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~42_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[3][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][10]~feeder .lut_mask = 16'hF0F0;
defparam \regs[3][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N11
dffeas \regs[3][10] (
	.clk(CLK),
	.d(\regs[3][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][10] .is_wysiwyg = "true";
defparam \regs[3][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N12
cycloneive_lcell_comb \Mux21~14 (
// Equation(s):
// \Mux21~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][10]~q ))) # (!dcifimemload_22 & (\regs[1][10]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[1][10]~q ),
	.datac(\regs[3][10]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux21~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~14 .lut_mask = 16'hA088;
defparam \Mux21~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N24
cycloneive_lcell_comb \Mux21~15 (
// Equation(s):
// \Mux21~15_combout  = (\Mux21~14_combout ) # ((\regs[2][10]~q  & (!dcifimemload_21 & dcifimemload_22)))

	.dataa(\regs[2][10]~q ),
	.datab(dcifimemload_21),
	.datac(\Mux21~14_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux21~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~15 .lut_mask = 16'hF2F0;
defparam \Mux21~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N18
cycloneive_lcell_comb \Mux21~16 (
// Equation(s):
// \Mux21~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux21~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & ((\Mux21~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux21~13_combout ),
	.datad(\Mux21~15_combout ),
	.cin(gnd),
	.combout(\Mux21~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~16 .lut_mask = 16'hB9A8;
defparam \Mux21~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y45_N16
cycloneive_lcell_comb \Mux21~19 (
// Equation(s):
// \Mux21~19_combout  = (dcifimemload_23 & ((\Mux21~16_combout  & ((\Mux21~18_combout ))) # (!\Mux21~16_combout  & (\Mux21~11_combout )))) # (!dcifimemload_23 & (((\Mux21~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux21~11_combout ),
	.datac(\Mux21~18_combout ),
	.datad(\Mux21~16_combout ),
	.cin(gnd),
	.combout(\Mux21~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~19 .lut_mask = 16'hF588;
defparam \Mux21~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N26
cycloneive_lcell_comb \regs~43 (
// Equation(s):
// \regs~43_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & ((ramiframload_9))) # (!cuifRegSel_0 & (Mux223))))

	.dataa(Mux221),
	.datab(cuifRegSel_11),
	.datac(ramiframload_9),
	.datad(cuifRegSel_0),
	.cin(gnd),
	.combout(\regs~43_combout ),
	.cout());
// synopsys translate_off
defparam \regs~43 .lut_mask = 16'h3022;
defparam \regs~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N14
cycloneive_lcell_comb \regs~44 (
// Equation(s):
// \regs~44_combout  = (!\Equal0~1_combout  & ((\regs~43_combout ) # ((\regs~64_combout  & \Add1~14_combout ))))

	.dataa(\Equal0~1_combout ),
	.datab(\regs~64_combout ),
	.datac(\regs~43_combout ),
	.datad(Add17),
	.cin(gnd),
	.combout(\regs~44_combout ),
	.cout());
// synopsys translate_off
defparam \regs~44 .lut_mask = 16'h5450;
defparam \regs~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N24
cycloneive_lcell_comb \regs[29][9]~feeder (
// Equation(s):
// \regs[29][9]~feeder_combout  = \regs~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[29][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][9]~feeder .lut_mask = 16'hF0F0;
defparam \regs[29][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N25
dffeas \regs[29][9] (
	.clk(CLK),
	.d(\regs[29][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][9] .is_wysiwyg = "true";
defparam \regs[29][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N16
cycloneive_lcell_comb \regs[21][9]~feeder (
// Equation(s):
// \regs[21][9]~feeder_combout  = \regs~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~44_combout ),
	.cin(gnd),
	.combout(\regs[21][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][9]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N17
dffeas \regs[21][9] (
	.clk(CLK),
	.d(\regs[21][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][9] .is_wysiwyg = "true";
defparam \regs[21][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N27
dffeas \regs[17][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][9] .is_wysiwyg = "true";
defparam \regs[17][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N9
dffeas \regs[25][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][9] .is_wysiwyg = "true";
defparam \regs[25][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N8
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[25][9]~q ))) # (!dcifimemload_19 & (\regs[17][9]~q ))))

	.dataa(dcifimemload_18),
	.datab(\regs[17][9]~q ),
	.datac(\regs[25][9]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hFA44;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N26
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (dcifimemload_18 & ((\Mux54~0_combout  & (\regs[29][9]~q )) # (!\Mux54~0_combout  & ((\regs[21][9]~q ))))) # (!dcifimemload_18 & (((\Mux54~0_combout ))))

	.dataa(\regs[29][9]~q ),
	.datab(\regs[21][9]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux54~0_combout ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hAFC0;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N25
dffeas \regs[24][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][9] .is_wysiwyg = "true";
defparam \regs[24][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N19
dffeas \regs[20][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][9] .is_wysiwyg = "true";
defparam \regs[20][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N18
cycloneive_lcell_comb \Mux54~4 (
// Equation(s):
// \Mux54~4_combout  = (dcifimemload_18 & (((\regs[20][9]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[16][9]~q  & ((!dcifimemload_19))))

	.dataa(\regs[16][9]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[20][9]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux54~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~4 .lut_mask = 16'hCCE2;
defparam \Mux54~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N24
cycloneive_lcell_comb \Mux54~5 (
// Equation(s):
// \Mux54~5_combout  = (dcifimemload_19 & ((\Mux54~4_combout  & (\regs[28][9]~q )) # (!\Mux54~4_combout  & ((\regs[24][9]~q ))))) # (!dcifimemload_19 & (((\Mux54~4_combout ))))

	.dataa(\regs[28][9]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[24][9]~q ),
	.datad(\Mux54~4_combout ),
	.cin(gnd),
	.combout(\Mux54~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~5 .lut_mask = 16'hBBC0;
defparam \Mux54~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N26
cycloneive_lcell_comb \regs[30][9]~feeder (
// Equation(s):
// \regs[30][9]~feeder_combout  = \regs~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~44_combout ),
	.cin(gnd),
	.combout(\regs[30][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[30][9]~feeder .lut_mask = 16'hFF00;
defparam \regs[30][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N27
dffeas \regs[30][9] (
	.clk(CLK),
	.d(\regs[30][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][9] .is_wysiwyg = "true";
defparam \regs[30][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N1
dffeas \regs[26][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][9] .is_wysiwyg = "true";
defparam \regs[26][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N23
dffeas \regs[18][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][9] .is_wysiwyg = "true";
defparam \regs[18][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N3
dffeas \regs[22][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][9] .is_wysiwyg = "true";
defparam \regs[22][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N2
cycloneive_lcell_comb \Mux54~2 (
// Equation(s):
// \Mux54~2_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\regs[22][9]~q ))) # (!dcifimemload_18 & (\regs[18][9]~q ))))

	.dataa(dcifimemload_19),
	.datab(\regs[18][9]~q ),
	.datac(\regs[22][9]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~2 .lut_mask = 16'hFA44;
defparam \Mux54~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N0
cycloneive_lcell_comb \Mux54~3 (
// Equation(s):
// \Mux54~3_combout  = (dcifimemload_19 & ((\Mux54~2_combout  & (\regs[30][9]~q )) # (!\Mux54~2_combout  & ((\regs[26][9]~q ))))) # (!dcifimemload_19 & (((\Mux54~2_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[30][9]~q ),
	.datac(\regs[26][9]~q ),
	.datad(\Mux54~2_combout ),
	.cin(gnd),
	.combout(\Mux54~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~3 .lut_mask = 16'hDDA0;
defparam \Mux54~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N4
cycloneive_lcell_comb \Mux54~6 (
// Equation(s):
// \Mux54~6_combout  = (dcifimemload_17 & (((dcifimemload_16) # (\Mux54~3_combout )))) # (!dcifimemload_17 & (\Mux54~5_combout  & (!dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\Mux54~5_combout ),
	.datac(dcifimemload_16),
	.datad(\Mux54~3_combout ),
	.cin(gnd),
	.combout(\Mux54~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~6 .lut_mask = 16'hAEA4;
defparam \Mux54~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N11
dffeas \regs[31][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][9] .is_wysiwyg = "true";
defparam \regs[31][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N3
dffeas \regs[23][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][9] .is_wysiwyg = "true";
defparam \regs[23][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N14
cycloneive_lcell_comb \regs[27][9]~feeder (
// Equation(s):
// \regs[27][9]~feeder_combout  = \regs~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~44_combout ),
	.cin(gnd),
	.combout(\regs[27][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][9]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N15
dffeas \regs[27][9] (
	.clk(CLK),
	.d(\regs[27][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][9] .is_wysiwyg = "true";
defparam \regs[27][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N8
cycloneive_lcell_comb \Mux54~7 (
// Equation(s):
// \Mux54~7_combout  = (dcifimemload_19 & (((\regs[27][9]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\regs[19][9]~q  & ((!dcifimemload_18))))

	.dataa(\regs[19][9]~q ),
	.datab(\regs[27][9]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux54~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~7 .lut_mask = 16'hF0CA;
defparam \Mux54~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N2
cycloneive_lcell_comb \Mux54~8 (
// Equation(s):
// \Mux54~8_combout  = (dcifimemload_18 & ((\Mux54~7_combout  & (\regs[31][9]~q )) # (!\Mux54~7_combout  & ((\regs[23][9]~q ))))) # (!dcifimemload_18 & (((\Mux54~7_combout ))))

	.dataa(\regs[31][9]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[23][9]~q ),
	.datad(\Mux54~7_combout ),
	.cin(gnd),
	.combout(\Mux54~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~8 .lut_mask = 16'hBBC0;
defparam \Mux54~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N15
dffeas \regs[15][9] (
	.clk(CLK),
	.d(\regs~44_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][9] .is_wysiwyg = "true";
defparam \regs[15][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N4
cycloneive_lcell_comb \regs[14][9]~feeder (
// Equation(s):
// \regs[14][9]~feeder_combout  = \regs~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~44_combout ),
	.cin(gnd),
	.combout(\regs[14][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][9]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N5
dffeas \regs[14][9] (
	.clk(CLK),
	.d(\regs[14][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][9] .is_wysiwyg = "true";
defparam \regs[14][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N1
dffeas \regs[13][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][9] .is_wysiwyg = "true";
defparam \regs[13][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N23
dffeas \regs[12][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][9] .is_wysiwyg = "true";
defparam \regs[12][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N22
cycloneive_lcell_comb \Mux54~17 (
// Equation(s):
// \Mux54~17_combout  = (dcifimemload_16 & ((\regs[13][9]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[12][9]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[13][9]~q ),
	.datac(\regs[12][9]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux54~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~17 .lut_mask = 16'hAAD8;
defparam \Mux54~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N30
cycloneive_lcell_comb \Mux54~18 (
// Equation(s):
// \Mux54~18_combout  = (\Mux54~17_combout  & ((\regs[15][9]~q ) # ((!dcifimemload_17)))) # (!\Mux54~17_combout  & (((\regs[14][9]~q  & dcifimemload_17))))

	.dataa(\regs[15][9]~q ),
	.datab(\regs[14][9]~q ),
	.datac(\Mux54~17_combout ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux54~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~18 .lut_mask = 16'hACF0;
defparam \Mux54~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N11
dffeas \regs[5][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][9] .is_wysiwyg = "true";
defparam \regs[5][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N10
cycloneive_lcell_comb \Mux54~10 (
// Equation(s):
// \Mux54~10_combout  = (dcifimemload_16 & (((\regs[5][9]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][9]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][9]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[5][9]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux54~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~10 .lut_mask = 16'hCCE2;
defparam \Mux54~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N19
dffeas \regs[7][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][9] .is_wysiwyg = "true";
defparam \regs[7][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N25
dffeas \regs[6][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][9] .is_wysiwyg = "true";
defparam \regs[6][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N24
cycloneive_lcell_comb \Mux54~11 (
// Equation(s):
// \Mux54~11_combout  = (\Mux54~10_combout  & ((\regs[7][9]~q ) # ((!dcifimemload_17)))) # (!\Mux54~10_combout  & (((\regs[6][9]~q  & dcifimemload_17))))

	.dataa(\Mux54~10_combout ),
	.datab(\regs[7][9]~q ),
	.datac(\regs[6][9]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux54~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~11 .lut_mask = 16'hD8AA;
defparam \Mux54~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N23
dffeas \regs[9][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][9] .is_wysiwyg = "true";
defparam \regs[9][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N31
dffeas \regs[11][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][9] .is_wysiwyg = "true";
defparam \regs[11][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N13
dffeas \regs[10][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][9] .is_wysiwyg = "true";
defparam \regs[10][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N29
dffeas \regs[8][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][9] .is_wysiwyg = "true";
defparam \regs[8][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N28
cycloneive_lcell_comb \Mux54~12 (
// Equation(s):
// \Mux54~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][9]~q )) # (!dcifimemload_17 & ((\regs[8][9]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][9]~q ),
	.datac(\regs[8][9]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux54~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~12 .lut_mask = 16'hEE50;
defparam \Mux54~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N30
cycloneive_lcell_comb \Mux54~13 (
// Equation(s):
// \Mux54~13_combout  = (dcifimemload_16 & ((\Mux54~12_combout  & ((\regs[11][9]~q ))) # (!\Mux54~12_combout  & (\regs[9][9]~q )))) # (!dcifimemload_16 & (((\Mux54~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][9]~q ),
	.datac(\regs[11][9]~q ),
	.datad(\Mux54~12_combout ),
	.cin(gnd),
	.combout(\Mux54~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~13 .lut_mask = 16'hF588;
defparam \Mux54~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y45_N1
dffeas \regs[2][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][9] .is_wysiwyg = "true";
defparam \regs[2][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y45_N19
dffeas \regs[1][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][9] .is_wysiwyg = "true";
defparam \regs[1][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N18
cycloneive_lcell_comb \Mux54~14 (
// Equation(s):
// \Mux54~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][9]~q )) # (!dcifimemload_17 & ((\regs[1][9]~q )))))

	.dataa(\regs[3][9]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][9]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux54~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~14 .lut_mask = 16'h88C0;
defparam \Mux54~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N0
cycloneive_lcell_comb \Mux54~15 (
// Equation(s):
// \Mux54~15_combout  = (\Mux54~14_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][9]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[2][9]~q ),
	.datad(\Mux54~14_combout ),
	.cin(gnd),
	.combout(\Mux54~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~15 .lut_mask = 16'hFF20;
defparam \Mux54~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N20
cycloneive_lcell_comb \Mux54~16 (
// Equation(s):
// \Mux54~16_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\Mux54~13_combout )) # (!dcifimemload_19 & ((\Mux54~15_combout )))))

	.dataa(\Mux54~13_combout ),
	.datab(dcifimemload_18),
	.datac(dcifimemload_19),
	.datad(\Mux54~15_combout ),
	.cin(gnd),
	.combout(\Mux54~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~16 .lut_mask = 16'hE3E0;
defparam \Mux54~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N13
dffeas \regs[19][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][9] .is_wysiwyg = "true";
defparam \regs[19][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N12
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// \Mux22~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[23][9]~q )) # (!dcifimemload_23 & ((\regs[19][9]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[23][9]~q ),
	.datac(\regs[19][9]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hEE50;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N10
cycloneive_lcell_comb \Mux22~8 (
// Equation(s):
// \Mux22~8_combout  = (dcifimemload_24 & ((\Mux22~7_combout  & ((\regs[31][9]~q ))) # (!\Mux22~7_combout  & (\regs[27][9]~q )))) # (!dcifimemload_24 & (((\Mux22~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][9]~q ),
	.datac(\regs[31][9]~q ),
	.datad(\Mux22~7_combout ),
	.cin(gnd),
	.combout(\Mux22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~8 .lut_mask = 16'hF588;
defparam \Mux22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N26
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[21][9]~q )) # (!dcifimemload_23 & ((\regs[17][9]~q )))))

	.dataa(\regs[21][9]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[17][9]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hEE30;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N8
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (dcifimemload_24 & ((\Mux22~0_combout  & ((\regs[29][9]~q ))) # (!\Mux22~0_combout  & (\regs[25][9]~q )))) # (!dcifimemload_24 & (((\Mux22~0_combout ))))

	.dataa(\regs[25][9]~q ),
	.datab(\regs[29][9]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hCFA0;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N16
cycloneive_lcell_comb \regs[16][9]~feeder (
// Equation(s):
// \regs[16][9]~feeder_combout  = \regs~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[16][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[16][9]~feeder .lut_mask = 16'hF0F0;
defparam \regs[16][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y45_N17
dffeas \regs[16][9] (
	.clk(CLK),
	.d(\regs[16][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][9] .is_wysiwyg = "true";
defparam \regs[16][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N4
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (dcifimemload_24 & (((\regs[24][9]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[16][9]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[16][9]~q ),
	.datac(\regs[24][9]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hAAE4;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N30
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// \Mux22~5_combout  = (\Mux22~4_combout  & ((\regs[28][9]~q ) # ((!dcifimemload_23)))) # (!\Mux22~4_combout  & (((\regs[20][9]~q  & dcifimemload_23))))

	.dataa(\regs[28][9]~q ),
	.datab(\regs[20][9]~q ),
	.datac(\Mux22~4_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hACF0;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N22
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (dcifimemload_24 & ((\regs[26][9]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[18][9]~q  & !dcifimemload_23))))

	.dataa(\regs[26][9]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[18][9]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hCCB8;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N6
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (\Mux22~2_combout  & ((\regs[30][9]~q ) # ((!dcifimemload_23)))) # (!\Mux22~2_combout  & (((\regs[22][9]~q  & dcifimemload_23))))

	.dataa(\regs[30][9]~q ),
	.datab(\Mux22~2_combout ),
	.datac(\regs[22][9]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hB8CC;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N2
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux22~3_combout ))) # (!dcifimemload_22 & (\Mux22~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux22~5_combout ),
	.datad(\Mux22~3_combout ),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hDC98;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N8
cycloneive_lcell_comb \Mux22~9 (
// Equation(s):
// \Mux22~9_combout  = (dcifimemload_21 & ((\Mux22~6_combout  & (\Mux22~8_combout )) # (!\Mux22~6_combout  & ((\Mux22~1_combout ))))) # (!dcifimemload_21 & (((\Mux22~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux22~8_combout ),
	.datac(\Mux22~1_combout ),
	.datad(\Mux22~6_combout ),
	.cin(gnd),
	.combout(\Mux22~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~9 .lut_mask = 16'hDDA0;
defparam \Mux22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N22
cycloneive_lcell_comb \Mux22~11 (
// Equation(s):
// \Mux22~11_combout  = (\Mux22~10_combout  & (((\regs[11][9]~q )) # (!dcifimemload_21))) # (!\Mux22~10_combout  & (dcifimemload_21 & (\regs[9][9]~q )))

	.dataa(\Mux22~10_combout ),
	.datab(dcifimemload_21),
	.datac(\regs[9][9]~q ),
	.datad(\regs[11][9]~q ),
	.cin(gnd),
	.combout(\Mux22~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~11 .lut_mask = 16'hEA62;
defparam \Mux22~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N0
cycloneive_lcell_comb \Mux22~17 (
// Equation(s):
// \Mux22~17_combout  = (dcifimemload_21 & (((\regs[13][9]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][9]~q  & ((!dcifimemload_22))))

	.dataa(\regs[12][9]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[13][9]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux22~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~17 .lut_mask = 16'hCCE2;
defparam \Mux22~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N14
cycloneive_lcell_comb \Mux22~18 (
// Equation(s):
// \Mux22~18_combout  = (dcifimemload_22 & ((\Mux22~17_combout  & (\regs[15][9]~q )) # (!\Mux22~17_combout  & ((\regs[14][9]~q ))))) # (!dcifimemload_22 & (((\Mux22~17_combout ))))

	.dataa(\regs[15][9]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[14][9]~q ),
	.datad(\Mux22~17_combout ),
	.cin(gnd),
	.combout(\Mux22~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~18 .lut_mask = 16'hBBC0;
defparam \Mux22~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N16
cycloneive_lcell_comb \regs[3][9]~feeder (
// Equation(s):
// \regs[3][9]~feeder_combout  = \regs~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[3][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][9]~feeder .lut_mask = 16'hF0F0;
defparam \regs[3][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N17
dffeas \regs[3][9] (
	.clk(CLK),
	.d(\regs[3][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][9] .is_wysiwyg = "true";
defparam \regs[3][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N0
cycloneive_lcell_comb \Mux22~14 (
// Equation(s):
// \Mux22~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\regs[3][9]~q )) # (!dcifimemload_22 & ((\regs[1][9]~q )))))

	.dataa(dcifimemload_21),
	.datab(\regs[3][9]~q ),
	.datac(dcifimemload_22),
	.datad(\regs[1][9]~q ),
	.cin(gnd),
	.combout(\Mux22~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~14 .lut_mask = 16'h8A80;
defparam \Mux22~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N26
cycloneive_lcell_comb \Mux22~15 (
// Equation(s):
// \Mux22~15_combout  = (\Mux22~14_combout ) # ((!dcifimemload_21 & (\regs[2][9]~q  & dcifimemload_22)))

	.dataa(dcifimemload_21),
	.datab(\regs[2][9]~q ),
	.datac(\Mux22~14_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux22~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~15 .lut_mask = 16'hF4F0;
defparam \Mux22~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N9
dffeas \regs[4][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~44_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][9] .is_wysiwyg = "true";
defparam \regs[4][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N8
cycloneive_lcell_comb \Mux22~12 (
// Equation(s):
// \Mux22~12_combout  = (dcifimemload_21 & ((dcifimemload_22) # ((\regs[5][9]~q )))) # (!dcifimemload_21 & (!dcifimemload_22 & (\regs[4][9]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[4][9]~q ),
	.datad(\regs[5][9]~q ),
	.cin(gnd),
	.combout(\Mux22~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~12 .lut_mask = 16'hBA98;
defparam \Mux22~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N18
cycloneive_lcell_comb \Mux22~13 (
// Equation(s):
// \Mux22~13_combout  = (dcifimemload_22 & ((\Mux22~12_combout  & ((\regs[7][9]~q ))) # (!\Mux22~12_combout  & (\regs[6][9]~q )))) # (!dcifimemload_22 & (((\Mux22~12_combout ))))

	.dataa(\regs[6][9]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[7][9]~q ),
	.datad(\Mux22~12_combout ),
	.cin(gnd),
	.combout(\Mux22~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~13 .lut_mask = 16'hF388;
defparam \Mux22~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N12
cycloneive_lcell_comb \Mux22~16 (
// Equation(s):
// \Mux22~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux22~13_combout ))) # (!dcifimemload_23 & (\Mux22~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux22~15_combout ),
	.datad(\Mux22~13_combout ),
	.cin(gnd),
	.combout(\Mux22~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~16 .lut_mask = 16'hDC98;
defparam \Mux22~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y45_N16
cycloneive_lcell_comb \Mux22~19 (
// Equation(s):
// \Mux22~19_combout  = (dcifimemload_24 & ((\Mux22~16_combout  & ((\Mux22~18_combout ))) # (!\Mux22~16_combout  & (\Mux22~11_combout )))) # (!dcifimemload_24 & (((\Mux22~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux22~11_combout ),
	.datac(\Mux22~18_combout ),
	.datad(\Mux22~16_combout ),
	.cin(gnd),
	.combout(\Mux22~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~19 .lut_mask = 16'hF588;
defparam \Mux22~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N12
cycloneive_lcell_comb \regs~45 (
// Equation(s):
// \regs~45_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & ((ramiframload_8))) # (!cuifRegSel_0 & (Mux233))))

	.dataa(Mux231),
	.datab(cuifRegSel_11),
	.datac(ramiframload_8),
	.datad(cuifRegSel_0),
	.cin(gnd),
	.combout(\regs~45_combout ),
	.cout());
// synopsys translate_off
defparam \regs~45 .lut_mask = 16'h3022;
defparam \regs~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N20
cycloneive_lcell_comb \regs~46 (
// Equation(s):
// \regs~46_combout  = (!\Equal0~1_combout  & ((\regs~45_combout ) # ((\regs~64_combout  & \Add1~12_combout ))))

	.dataa(\Equal0~1_combout ),
	.datab(\regs~64_combout ),
	.datac(Add16),
	.datad(\regs~45_combout ),
	.cin(gnd),
	.combout(\regs~46_combout ),
	.cout());
// synopsys translate_off
defparam \regs~46 .lut_mask = 16'h5540;
defparam \regs~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N17
dffeas \regs[22][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][8] .is_wysiwyg = "true";
defparam \regs[22][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N7
dffeas \regs[30][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][8] .is_wysiwyg = "true";
defparam \regs[30][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N16
cycloneive_lcell_comb \Mux55~3 (
// Equation(s):
// \Mux55~3_combout  = (\Mux55~2_combout  & (((\regs[30][8]~q )) # (!dcifimemload_18))) # (!\Mux55~2_combout  & (dcifimemload_18 & (\regs[22][8]~q )))

	.dataa(\Mux55~2_combout ),
	.datab(dcifimemload_18),
	.datac(\regs[22][8]~q ),
	.datad(\regs[30][8]~q ),
	.cin(gnd),
	.combout(\Mux55~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~3 .lut_mask = 16'hEA62;
defparam \Mux55~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N25
dffeas \regs[20][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][8] .is_wysiwyg = "true";
defparam \regs[20][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N7
dffeas \regs[24][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][8] .is_wysiwyg = "true";
defparam \regs[24][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N6
cycloneive_lcell_comb \Mux55~4 (
// Equation(s):
// \Mux55~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[24][8]~q ))) # (!dcifimemload_19 & (\regs[16][8]~q ))))

	.dataa(\regs[16][8]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[24][8]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux55~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~4 .lut_mask = 16'hFC22;
defparam \Mux55~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N24
cycloneive_lcell_comb \Mux55~5 (
// Equation(s):
// \Mux55~5_combout  = (dcifimemload_18 & ((\Mux55~4_combout  & (\regs[28][8]~q )) # (!\Mux55~4_combout  & ((\regs[20][8]~q ))))) # (!dcifimemload_18 & (((\Mux55~4_combout ))))

	.dataa(\regs[28][8]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[20][8]~q ),
	.datad(\Mux55~4_combout ),
	.cin(gnd),
	.combout(\Mux55~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~5 .lut_mask = 16'hBBC0;
defparam \Mux55~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N4
cycloneive_lcell_comb \Mux55~6 (
// Equation(s):
// \Mux55~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux55~3_combout )) # (!dcifimemload_17 & ((\Mux55~5_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux55~3_combout ),
	.datad(\Mux55~5_combout ),
	.cin(gnd),
	.combout(\Mux55~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~6 .lut_mask = 16'hD9C8;
defparam \Mux55~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N22
cycloneive_lcell_comb \regs[29][8]~feeder (
// Equation(s):
// \regs[29][8]~feeder_combout  = \regs~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~46_combout ),
	.cin(gnd),
	.combout(\regs[29][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][8]~feeder .lut_mask = 16'hFF00;
defparam \regs[29][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N23
dffeas \regs[29][8] (
	.clk(CLK),
	.d(\regs[29][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][8] .is_wysiwyg = "true";
defparam \regs[29][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N3
dffeas \regs[25][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][8] .is_wysiwyg = "true";
defparam \regs[25][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N29
dffeas \regs[17][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][8] .is_wysiwyg = "true";
defparam \regs[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N12
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[21][8]~q )) # (!dcifimemload_18 & ((\regs[17][8]~q )))))

	.dataa(\regs[21][8]~q ),
	.datab(\regs[17][8]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hFA0C;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N2
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (dcifimemload_19 & ((\Mux55~0_combout  & (\regs[29][8]~q )) # (!\Mux55~0_combout  & ((\regs[25][8]~q ))))) # (!dcifimemload_19 & (((\Mux55~0_combout ))))

	.dataa(\regs[29][8]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[25][8]~q ),
	.datad(\Mux55~0_combout ),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hBBC0;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N23
dffeas \regs[31][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][8] .is_wysiwyg = "true";
defparam \regs[31][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N23
dffeas \regs[27][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][8] .is_wysiwyg = "true";
defparam \regs[27][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N5
dffeas \regs[19][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][8] .is_wysiwyg = "true";
defparam \regs[19][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N2
cycloneive_lcell_comb \Mux55~7 (
// Equation(s):
// \Mux55~7_combout  = (dcifimemload_18 & ((\regs[23][8]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[19][8]~q  & !dcifimemload_19))))

	.dataa(\regs[23][8]~q ),
	.datab(\regs[19][8]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux55~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~7 .lut_mask = 16'hF0AC;
defparam \Mux55~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N22
cycloneive_lcell_comb \Mux55~8 (
// Equation(s):
// \Mux55~8_combout  = (dcifimemload_19 & ((\Mux55~7_combout  & (\regs[31][8]~q )) # (!\Mux55~7_combout  & ((\regs[27][8]~q ))))) # (!dcifimemload_19 & (((\Mux55~7_combout ))))

	.dataa(\regs[31][8]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[27][8]~q ),
	.datad(\Mux55~7_combout ),
	.cin(gnd),
	.combout(\Mux55~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~8 .lut_mask = 16'hBBC0;
defparam \Mux55~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N21
dffeas \regs[11][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][8] .is_wysiwyg = "true";
defparam \regs[11][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N25
dffeas \regs[9][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][8] .is_wysiwyg = "true";
defparam \regs[9][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N19
dffeas \regs[10][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][8] .is_wysiwyg = "true";
defparam \regs[10][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N18
cycloneive_lcell_comb \Mux55~10 (
// Equation(s):
// \Mux55~10_combout  = (dcifimemload_17 & (((\regs[10][8]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\regs[8][8]~q  & ((!dcifimemload_16))))

	.dataa(\regs[8][8]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[10][8]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux55~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~10 .lut_mask = 16'hCCE2;
defparam \Mux55~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N24
cycloneive_lcell_comb \Mux55~11 (
// Equation(s):
// \Mux55~11_combout  = (dcifimemload_16 & ((\Mux55~10_combout  & (\regs[11][8]~q )) # (!\Mux55~10_combout  & ((\regs[9][8]~q ))))) # (!dcifimemload_16 & (((\Mux55~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[11][8]~q ),
	.datac(\regs[9][8]~q ),
	.datad(\Mux55~10_combout ),
	.cin(gnd),
	.combout(\Mux55~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~11 .lut_mask = 16'hDDA0;
defparam \Mux55~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N21
dffeas \regs[15][8] (
	.clk(CLK),
	.d(\regs~46_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][8] .is_wysiwyg = "true";
defparam \regs[15][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y44_N25
dffeas \regs[14][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][8] .is_wysiwyg = "true";
defparam \regs[14][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y44_N19
dffeas \regs[12][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][8] .is_wysiwyg = "true";
defparam \regs[12][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N18
cycloneive_lcell_comb \Mux55~17 (
// Equation(s):
// \Mux55~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][8]~q )) # (!dcifimemload_16 & ((\regs[12][8]~q )))))

	.dataa(\regs[13][8]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][8]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux55~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~17 .lut_mask = 16'hEE30;
defparam \Mux55~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N24
cycloneive_lcell_comb \Mux55~18 (
// Equation(s):
// \Mux55~18_combout  = (dcifimemload_17 & ((\Mux55~17_combout  & (\regs[15][8]~q )) # (!\Mux55~17_combout  & ((\regs[14][8]~q ))))) # (!dcifimemload_17 & (((\Mux55~17_combout ))))

	.dataa(\regs[15][8]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[14][8]~q ),
	.datad(\Mux55~17_combout ),
	.cin(gnd),
	.combout(\Mux55~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~18 .lut_mask = 16'hBBC0;
defparam \Mux55~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y45_N21
dffeas \regs[2][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][8] .is_wysiwyg = "true";
defparam \regs[2][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N2
cycloneive_lcell_comb \regs[3][8]~feeder (
// Equation(s):
// \regs[3][8]~feeder_combout  = \regs~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~46_combout ),
	.cin(gnd),
	.combout(\regs[3][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][8]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N3
dffeas \regs[3][8] (
	.clk(CLK),
	.d(\regs[3][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][8] .is_wysiwyg = "true";
defparam \regs[3][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y45_N7
dffeas \regs[1][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][8] .is_wysiwyg = "true";
defparam \regs[1][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N6
cycloneive_lcell_comb \Mux55~14 (
// Equation(s):
// \Mux55~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][8]~q )) # (!dcifimemload_17 & ((\regs[1][8]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[3][8]~q ),
	.datac(\regs[1][8]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux55~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~14 .lut_mask = 16'h88A0;
defparam \Mux55~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N20
cycloneive_lcell_comb \Mux55~15 (
// Equation(s):
// \Mux55~15_combout  = (\Mux55~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][8]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][8]~q ),
	.datad(\Mux55~14_combout ),
	.cin(gnd),
	.combout(\Mux55~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~15 .lut_mask = 16'hFF40;
defparam \Mux55~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N3
dffeas \regs[6][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][8] .is_wysiwyg = "true";
defparam \regs[6][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N17
dffeas \regs[7][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][8] .is_wysiwyg = "true";
defparam \regs[7][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N27
dffeas \regs[5][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][8] .is_wysiwyg = "true";
defparam \regs[5][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N15
dffeas \regs[4][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][8] .is_wysiwyg = "true";
defparam \regs[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N14
cycloneive_lcell_comb \Mux55~12 (
// Equation(s):
// \Mux55~12_combout  = (dcifimemload_16 & ((\regs[5][8]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][8]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[5][8]~q ),
	.datac(\regs[4][8]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux55~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~12 .lut_mask = 16'hAAD8;
defparam \Mux55~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N16
cycloneive_lcell_comb \Mux55~13 (
// Equation(s):
// \Mux55~13_combout  = (dcifimemload_17 & ((\Mux55~12_combout  & ((\regs[7][8]~q ))) # (!\Mux55~12_combout  & (\regs[6][8]~q )))) # (!dcifimemload_17 & (((\Mux55~12_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][8]~q ),
	.datac(\regs[7][8]~q ),
	.datad(\Mux55~12_combout ),
	.cin(gnd),
	.combout(\Mux55~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~13 .lut_mask = 16'hF588;
defparam \Mux55~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N18
cycloneive_lcell_comb \Mux55~16 (
// Equation(s):
// \Mux55~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux55~13_combout ))) # (!dcifimemload_18 & (\Mux55~15_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux55~15_combout ),
	.datad(\Mux55~13_combout ),
	.cin(gnd),
	.combout(\Mux55~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~16 .lut_mask = 16'hDC98;
defparam \Mux55~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N29
dffeas \regs[18][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][8] .is_wysiwyg = "true";
defparam \regs[18][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N28
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (dcifimemload_23 & ((\regs[22][8]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[18][8]~q  & !dcifimemload_24))))

	.dataa(\regs[22][8]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[18][8]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hCCB8;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N6
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (\Mux23~2_combout  & (((\regs[30][8]~q ) # (!dcifimemload_24)))) # (!\Mux23~2_combout  & (\regs[26][8]~q  & ((dcifimemload_24))))

	.dataa(\regs[26][8]~q ),
	.datab(\Mux23~2_combout ),
	.datac(\regs[30][8]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hE2CC;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N21
dffeas \regs[28][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][8] .is_wysiwyg = "true";
defparam \regs[28][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y42_N11
dffeas \regs[16][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][8] .is_wysiwyg = "true";
defparam \regs[16][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N10
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (dcifimemload_23 & ((\regs[20][8]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[16][8]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[20][8]~q ),
	.datac(\regs[16][8]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hAAD8;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N20
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (dcifimemload_24 & ((\Mux23~4_combout  & ((\regs[28][8]~q ))) # (!\Mux23~4_combout  & (\regs[24][8]~q )))) # (!dcifimemload_24 & (((\Mux23~4_combout ))))

	.dataa(\regs[24][8]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[28][8]~q ),
	.datad(\Mux23~4_combout ),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hF388;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N26
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux23~3_combout )) # (!dcifimemload_22 & ((\Mux23~5_combout )))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux23~3_combout ),
	.datad(\Mux23~5_combout ),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hD9C8;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N20
cycloneive_lcell_comb \regs[21][8]~feeder (
// Equation(s):
// \regs[21][8]~feeder_combout  = \regs~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~46_combout ),
	.cin(gnd),
	.combout(\regs[21][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][8]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N21
dffeas \regs[21][8] (
	.clk(CLK),
	.d(\regs[21][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][8] .is_wysiwyg = "true";
defparam \regs[21][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N28
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (dcifimemload_24 & ((\regs[25][8]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[17][8]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[25][8]~q ),
	.datac(\regs[17][8]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hAAD8;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N8
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (dcifimemload_23 & ((\Mux23~0_combout  & (\regs[29][8]~q )) # (!\Mux23~0_combout  & ((\regs[21][8]~q ))))) # (!dcifimemload_23 & (((\Mux23~0_combout ))))

	.dataa(\regs[29][8]~q ),
	.datab(\regs[21][8]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux23~0_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hAFC0;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N4
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// \Mux23~7_combout  = (dcifimemload_24 & ((\regs[27][8]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[19][8]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[27][8]~q ),
	.datac(\regs[19][8]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hAAD8;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N22
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// \Mux23~8_combout  = (\Mux23~7_combout  & (((\regs[31][8]~q ) # (!dcifimemload_23)))) # (!\Mux23~7_combout  & (\regs[23][8]~q  & ((dcifimemload_23))))

	.dataa(\regs[23][8]~q ),
	.datab(\Mux23~7_combout ),
	.datac(\regs[31][8]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'hE2CC;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N16
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// \Mux23~9_combout  = (\Mux23~6_combout  & (((\Mux23~8_combout )) # (!dcifimemload_21))) # (!\Mux23~6_combout  & (dcifimemload_21 & (\Mux23~1_combout )))

	.dataa(\Mux23~6_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux23~1_combout ),
	.datad(\Mux23~8_combout ),
	.cin(gnd),
	.combout(\Mux23~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hEA62;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N16
cycloneive_lcell_comb \regs[13][8]~feeder (
// Equation(s):
// \regs[13][8]~feeder_combout  = \regs~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~46_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[13][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][8]~feeder .lut_mask = 16'hF0F0;
defparam \regs[13][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y44_N17
dffeas \regs[13][8] (
	.clk(CLK),
	.d(\regs[13][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][8] .is_wysiwyg = "true";
defparam \regs[13][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N22
cycloneive_lcell_comb \Mux23~17 (
// Equation(s):
// \Mux23~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\regs[13][8]~q ))) # (!dcifimemload_21 & (\regs[12][8]~q ))))

	.dataa(dcifimemload_22),
	.datab(\regs[12][8]~q ),
	.datac(\regs[13][8]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux23~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~17 .lut_mask = 16'hFA44;
defparam \Mux23~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N22
cycloneive_lcell_comb \Mux23~18 (
// Equation(s):
// \Mux23~18_combout  = (dcifimemload_22 & ((\Mux23~17_combout  & ((\regs[15][8]~q ))) # (!\Mux23~17_combout  & (\regs[14][8]~q )))) # (!dcifimemload_22 & (((\Mux23~17_combout ))))

	.dataa(\regs[14][8]~q ),
	.datab(dcifimemload_22),
	.datac(\Mux23~17_combout ),
	.datad(\regs[15][8]~q ),
	.cin(gnd),
	.combout(\Mux23~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~18 .lut_mask = 16'hF838;
defparam \Mux23~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N26
cycloneive_lcell_comb \Mux23~10 (
// Equation(s):
// \Mux23~10_combout  = (dcifimemload_21 & (((\regs[5][8]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][8]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][8]~q ),
	.datac(\regs[5][8]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux23~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~10 .lut_mask = 16'hAAE4;
defparam \Mux23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N2
cycloneive_lcell_comb \Mux23~11 (
// Equation(s):
// \Mux23~11_combout  = (dcifimemload_22 & ((\Mux23~10_combout  & (\regs[7][8]~q )) # (!\Mux23~10_combout  & ((\regs[6][8]~q ))))) # (!dcifimemload_22 & (((\Mux23~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[7][8]~q ),
	.datac(\regs[6][8]~q ),
	.datad(\Mux23~10_combout ),
	.cin(gnd),
	.combout(\Mux23~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~11 .lut_mask = 16'hDDA0;
defparam \Mux23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N11
dffeas \regs[8][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~46_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][8] .is_wysiwyg = "true";
defparam \regs[8][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N10
cycloneive_lcell_comb \Mux23~12 (
// Equation(s):
// \Mux23~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\regs[10][8]~q )) # (!dcifimemload_22 & ((\regs[8][8]~q )))))

	.dataa(\regs[10][8]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[8][8]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux23~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~12 .lut_mask = 16'hEE30;
defparam \Mux23~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N20
cycloneive_lcell_comb \Mux23~13 (
// Equation(s):
// \Mux23~13_combout  = (dcifimemload_21 & ((\Mux23~12_combout  & ((\regs[11][8]~q ))) # (!\Mux23~12_combout  & (\regs[9][8]~q )))) # (!dcifimemload_21 & (((\Mux23~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\regs[9][8]~q ),
	.datac(\regs[11][8]~q ),
	.datad(\Mux23~12_combout ),
	.cin(gnd),
	.combout(\Mux23~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~13 .lut_mask = 16'hF588;
defparam \Mux23~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N18
cycloneive_lcell_comb \Mux23~14 (
// Equation(s):
// \Mux23~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][8]~q ))) # (!dcifimemload_22 & (\regs[1][8]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[1][8]~q ),
	.datac(dcifimemload_22),
	.datad(\regs[3][8]~q ),
	.cin(gnd),
	.combout(\Mux23~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~14 .lut_mask = 16'hA808;
defparam \Mux23~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N2
cycloneive_lcell_comb \Mux23~15 (
// Equation(s):
// \Mux23~15_combout  = (\Mux23~14_combout ) # ((dcifimemload_22 & (\regs[2][8]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\regs[2][8]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux23~14_combout ),
	.cin(gnd),
	.combout(\Mux23~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~15 .lut_mask = 16'hFF08;
defparam \Mux23~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N0
cycloneive_lcell_comb \Mux23~16 (
// Equation(s):
// \Mux23~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux23~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & ((\Mux23~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux23~13_combout ),
	.datad(\Mux23~15_combout ),
	.cin(gnd),
	.combout(\Mux23~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~16 .lut_mask = 16'hB9A8;
defparam \Mux23~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y45_N12
cycloneive_lcell_comb \Mux23~19 (
// Equation(s):
// \Mux23~19_combout  = (dcifimemload_23 & ((\Mux23~16_combout  & (\Mux23~18_combout )) # (!\Mux23~16_combout  & ((\Mux23~11_combout ))))) # (!dcifimemload_23 & (((\Mux23~16_combout ))))

	.dataa(\Mux23~18_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux23~11_combout ),
	.datad(\Mux23~16_combout ),
	.cin(gnd),
	.combout(\Mux23~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~19 .lut_mask = 16'hBBC0;
defparam \Mux23~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N18
cycloneive_lcell_comb \regs~47 (
// Equation(s):
// \regs~47_combout  = (\Add1~10_combout  & (cuifRegSel_11 & !cuifRegSel_0))

	.dataa(Add15),
	.datab(cuifRegSel_11),
	.datac(gnd),
	.datad(cuifRegSel_0),
	.cin(gnd),
	.combout(\regs~47_combout ),
	.cout());
// synopsys translate_off
defparam \regs~47 .lut_mask = 16'h0088;
defparam \regs~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N4
cycloneive_lcell_comb \regs~48 (
// Equation(s):
// \regs~48_combout  = (cuifRegSel_0 & (ramiframload_7)) # (!cuifRegSel_0 & (((Mux241 & !Selector0))))

	.dataa(cuifRegSel_0),
	.datab(ramiframload_7),
	.datac(Mux241),
	.datad(Selector0),
	.cin(gnd),
	.combout(\regs~48_combout ),
	.cout());
// synopsys translate_off
defparam \regs~48 .lut_mask = 16'h88D8;
defparam \regs~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N14
cycloneive_lcell_comb \regs~49 (
// Equation(s):
// \regs~49_combout  = (!\Equal0~1_combout  & ((\regs~47_combout ) # ((!cuifRegSel_11 & \regs~48_combout ))))

	.dataa(cuifRegSel_11),
	.datab(\regs~47_combout ),
	.datac(\regs~48_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\regs~49_combout ),
	.cout());
// synopsys translate_off
defparam \regs~49 .lut_mask = 16'h00DC;
defparam \regs~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N15
dffeas \regs[21][7] (
	.clk(CLK),
	.d(\regs~49_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][7] .is_wysiwyg = "true";
defparam \regs[21][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N21
dffeas \regs[29][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][7] .is_wysiwyg = "true";
defparam \regs[29][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N11
dffeas \regs[17][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][7] .is_wysiwyg = "true";
defparam \regs[17][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N3
dffeas \regs[25][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][7] .is_wysiwyg = "true";
defparam \regs[25][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N2
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[25][7]~q ))) # (!dcifimemload_19 & (\regs[17][7]~q ))))

	.dataa(dcifimemload_18),
	.datab(\regs[17][7]~q ),
	.datac(\regs[25][7]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hFA44;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N22
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (dcifimemload_18 & ((\Mux56~0_combout  & ((\regs[29][7]~q ))) # (!\Mux56~0_combout  & (\regs[21][7]~q )))) # (!dcifimemload_18 & (((\Mux56~0_combout ))))

	.dataa(\regs[21][7]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[29][7]~q ),
	.datad(\Mux56~0_combout ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hF388;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N24
cycloneive_lcell_comb \regs[30][7]~feeder (
// Equation(s):
// \regs[30][7]~feeder_combout  = \regs~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~49_combout ),
	.cin(gnd),
	.combout(\regs[30][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[30][7]~feeder .lut_mask = 16'hFF00;
defparam \regs[30][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y45_N25
dffeas \regs[30][7] (
	.clk(CLK),
	.d(\regs[30][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][7] .is_wysiwyg = "true";
defparam \regs[30][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N13
dffeas \regs[26][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][7] .is_wysiwyg = "true";
defparam \regs[26][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N12
cycloneive_lcell_comb \Mux56~3 (
// Equation(s):
// \Mux56~3_combout  = (\Mux56~2_combout  & ((\regs[30][7]~q ) # ((!dcifimemload_19)))) # (!\Mux56~2_combout  & (((\regs[26][7]~q  & dcifimemload_19))))

	.dataa(\Mux56~2_combout ),
	.datab(\regs[30][7]~q ),
	.datac(\regs[26][7]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~3 .lut_mask = 16'hD8AA;
defparam \Mux56~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N25
dffeas \regs[24][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][7] .is_wysiwyg = "true";
defparam \regs[24][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N31
dffeas \regs[20][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][7] .is_wysiwyg = "true";
defparam \regs[20][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N30
cycloneive_lcell_comb \Mux56~4 (
// Equation(s):
// \Mux56~4_combout  = (dcifimemload_18 & (((\regs[20][7]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[16][7]~q  & ((!dcifimemload_19))))

	.dataa(\regs[16][7]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[20][7]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~4 .lut_mask = 16'hCCE2;
defparam \Mux56~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N24
cycloneive_lcell_comb \Mux56~5 (
// Equation(s):
// \Mux56~5_combout  = (dcifimemload_19 & ((\Mux56~4_combout  & (\regs[28][7]~q )) # (!\Mux56~4_combout  & ((\regs[24][7]~q ))))) # (!dcifimemload_19 & (((\Mux56~4_combout ))))

	.dataa(\regs[28][7]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[24][7]~q ),
	.datad(\Mux56~4_combout ),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~5 .lut_mask = 16'hBBC0;
defparam \Mux56~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N8
cycloneive_lcell_comb \Mux56~6 (
// Equation(s):
// \Mux56~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux56~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & ((\Mux56~5_combout ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux56~3_combout ),
	.datad(\Mux56~5_combout ),
	.cin(gnd),
	.combout(\Mux56~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~6 .lut_mask = 16'hB9A8;
defparam \Mux56~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N31
dffeas \regs[31][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][7] .is_wysiwyg = "true";
defparam \regs[31][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N19
dffeas \regs[23][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][7] .is_wysiwyg = "true";
defparam \regs[23][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N0
cycloneive_lcell_comb \regs[19][7]~feeder (
// Equation(s):
// \regs[19][7]~feeder_combout  = \regs~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~49_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[19][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][7]~feeder .lut_mask = 16'hF0F0;
defparam \regs[19][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N1
dffeas \regs[19][7] (
	.clk(CLK),
	.d(\regs[19][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][7] .is_wysiwyg = "true";
defparam \regs[19][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N19
dffeas \regs[27][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][7] .is_wysiwyg = "true";
defparam \regs[27][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N18
cycloneive_lcell_comb \Mux56~7 (
// Equation(s):
// \Mux56~7_combout  = (dcifimemload_19 & (((\regs[27][7]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\regs[19][7]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\regs[19][7]~q ),
	.datac(\regs[27][7]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux56~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~7 .lut_mask = 16'hAAE4;
defparam \Mux56~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N18
cycloneive_lcell_comb \Mux56~8 (
// Equation(s):
// \Mux56~8_combout  = (dcifimemload_18 & ((\Mux56~7_combout  & (\regs[31][7]~q )) # (!\Mux56~7_combout  & ((\regs[23][7]~q ))))) # (!dcifimemload_18 & (((\Mux56~7_combout ))))

	.dataa(\regs[31][7]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[23][7]~q ),
	.datad(\Mux56~7_combout ),
	.cin(gnd),
	.combout(\Mux56~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~8 .lut_mask = 16'hBBC0;
defparam \Mux56~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y44_N11
dffeas \regs[14][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][7] .is_wysiwyg = "true";
defparam \regs[14][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y44_N5
dffeas \regs[15][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][7] .is_wysiwyg = "true";
defparam \regs[15][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N16
cycloneive_lcell_comb \regs[13][7]~feeder (
// Equation(s):
// \regs[13][7]~feeder_combout  = \regs~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~49_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[13][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][7]~feeder .lut_mask = 16'hF0F0;
defparam \regs[13][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N17
dffeas \regs[13][7] (
	.clk(CLK),
	.d(\regs[13][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][7] .is_wysiwyg = "true";
defparam \regs[13][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N19
dffeas \regs[12][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][7] .is_wysiwyg = "true";
defparam \regs[12][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N18
cycloneive_lcell_comb \Mux56~17 (
// Equation(s):
// \Mux56~17_combout  = (dcifimemload_16 & ((\regs[13][7]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[12][7]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[13][7]~q ),
	.datac(\regs[12][7]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux56~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~17 .lut_mask = 16'hAAD8;
defparam \Mux56~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N4
cycloneive_lcell_comb \Mux56~18 (
// Equation(s):
// \Mux56~18_combout  = (dcifimemload_17 & ((\Mux56~17_combout  & ((\regs[15][7]~q ))) # (!\Mux56~17_combout  & (\regs[14][7]~q )))) # (!dcifimemload_17 & (((\Mux56~17_combout ))))

	.dataa(\regs[14][7]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[15][7]~q ),
	.datad(\Mux56~17_combout ),
	.cin(gnd),
	.combout(\Mux56~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~18 .lut_mask = 16'hF388;
defparam \Mux56~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N11
dffeas \regs[7][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][7] .is_wysiwyg = "true";
defparam \regs[7][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N13
dffeas \regs[6][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][7] .is_wysiwyg = "true";
defparam \regs[6][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N3
dffeas \regs[5][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][7] .is_wysiwyg = "true";
defparam \regs[5][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N2
cycloneive_lcell_comb \Mux56~10 (
// Equation(s):
// \Mux56~10_combout  = (dcifimemload_16 & (((\regs[5][7]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][7]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][7]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[5][7]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux56~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~10 .lut_mask = 16'hCCE2;
defparam \Mux56~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N12
cycloneive_lcell_comb \Mux56~11 (
// Equation(s):
// \Mux56~11_combout  = (dcifimemload_17 & ((\Mux56~10_combout  & (\regs[7][7]~q )) # (!\Mux56~10_combout  & ((\regs[6][7]~q ))))) # (!dcifimemload_17 & (((\Mux56~10_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[7][7]~q ),
	.datac(\regs[6][7]~q ),
	.datad(\Mux56~10_combout ),
	.cin(gnd),
	.combout(\Mux56~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~11 .lut_mask = 16'hDDA0;
defparam \Mux56~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N17
dffeas \regs[10][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][7] .is_wysiwyg = "true";
defparam \regs[10][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N9
dffeas \regs[8][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][7] .is_wysiwyg = "true";
defparam \regs[8][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N8
cycloneive_lcell_comb \Mux56~12 (
// Equation(s):
// \Mux56~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][7]~q )) # (!dcifimemload_17 & ((\regs[8][7]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][7]~q ),
	.datac(\regs[8][7]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux56~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~12 .lut_mask = 16'hEE50;
defparam \Mux56~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N11
dffeas \regs[11][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][7] .is_wysiwyg = "true";
defparam \regs[11][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N7
dffeas \regs[9][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][7] .is_wysiwyg = "true";
defparam \regs[9][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N10
cycloneive_lcell_comb \Mux56~13 (
// Equation(s):
// \Mux56~13_combout  = (dcifimemload_16 & ((\Mux56~12_combout  & (\regs[11][7]~q )) # (!\Mux56~12_combout  & ((\regs[9][7]~q ))))) # (!dcifimemload_16 & (\Mux56~12_combout ))

	.dataa(dcifimemload_16),
	.datab(\Mux56~12_combout ),
	.datac(\regs[11][7]~q ),
	.datad(\regs[9][7]~q ),
	.cin(gnd),
	.combout(\Mux56~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~13 .lut_mask = 16'hE6C4;
defparam \Mux56~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y45_N23
dffeas \regs[2][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][7] .is_wysiwyg = "true";
defparam \regs[2][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y45_N1
dffeas \regs[1][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][7] .is_wysiwyg = "true";
defparam \regs[1][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N0
cycloneive_lcell_comb \Mux56~14 (
// Equation(s):
// \Mux56~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][7]~q )) # (!dcifimemload_17 & ((\regs[1][7]~q )))))

	.dataa(\regs[3][7]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][7]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux56~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~14 .lut_mask = 16'h88C0;
defparam \Mux56~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N22
cycloneive_lcell_comb \Mux56~15 (
// Equation(s):
// \Mux56~15_combout  = (\Mux56~14_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][7]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[2][7]~q ),
	.datad(\Mux56~14_combout ),
	.cin(gnd),
	.combout(\Mux56~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~15 .lut_mask = 16'hFF20;
defparam \Mux56~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N28
cycloneive_lcell_comb \Mux56~16 (
// Equation(s):
// \Mux56~16_combout  = (dcifimemload_19 & ((\Mux56~13_combout ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((!dcifimemload_18 & \Mux56~15_combout ))))

	.dataa(\Mux56~13_combout ),
	.datab(dcifimemload_19),
	.datac(dcifimemload_18),
	.datad(\Mux56~15_combout ),
	.cin(gnd),
	.combout(\Mux56~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~16 .lut_mask = 16'hCBC8;
defparam \Mux56~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N16
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][7]~q ))) # (!dcifimemload_22 & (\regs[8][7]~q ))))

	.dataa(\regs[8][7]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[10][7]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'hFC22;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N6
cycloneive_lcell_comb \Mux24~11 (
// Equation(s):
// \Mux24~11_combout  = (dcifimemload_21 & ((\Mux24~10_combout  & (\regs[11][7]~q )) # (!\Mux24~10_combout  & ((\regs[9][7]~q ))))) # (!dcifimemload_21 & (((\Mux24~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\regs[11][7]~q ),
	.datac(\regs[9][7]~q ),
	.datad(\Mux24~10_combout ),
	.cin(gnd),
	.combout(\Mux24~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~11 .lut_mask = 16'hDDA0;
defparam \Mux24~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N18
cycloneive_lcell_comb \Mux24~17 (
// Equation(s):
// \Mux24~17_combout  = (dcifimemload_21 & (((\regs[13][7]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][7]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][7]~q ),
	.datac(\regs[13][7]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux24~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~17 .lut_mask = 16'hAAE4;
defparam \Mux24~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y44_N10
cycloneive_lcell_comb \Mux24~18 (
// Equation(s):
// \Mux24~18_combout  = (dcifimemload_22 & ((\Mux24~17_combout  & (\regs[15][7]~q )) # (!\Mux24~17_combout  & ((\regs[14][7]~q ))))) # (!dcifimemload_22 & (((\Mux24~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][7]~q ),
	.datac(\regs[14][7]~q ),
	.datad(\Mux24~17_combout ),
	.cin(gnd),
	.combout(\Mux24~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~18 .lut_mask = 16'hDDA0;
defparam \Mux24~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N21
dffeas \regs[4][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][7] .is_wysiwyg = "true";
defparam \regs[4][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N20
cycloneive_lcell_comb \Mux24~12 (
// Equation(s):
// \Mux24~12_combout  = (dcifimemload_21 & ((dcifimemload_22) # ((\regs[5][7]~q )))) # (!dcifimemload_21 & (!dcifimemload_22 & (\regs[4][7]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[4][7]~q ),
	.datad(\regs[5][7]~q ),
	.cin(gnd),
	.combout(\Mux24~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~12 .lut_mask = 16'hBA98;
defparam \Mux24~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N10
cycloneive_lcell_comb \Mux24~13 (
// Equation(s):
// \Mux24~13_combout  = (dcifimemload_22 & ((\Mux24~12_combout  & ((\regs[7][7]~q ))) # (!\Mux24~12_combout  & (\regs[6][7]~q )))) # (!dcifimemload_22 & (((\Mux24~12_combout ))))

	.dataa(\regs[6][7]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[7][7]~q ),
	.datad(\Mux24~12_combout ),
	.cin(gnd),
	.combout(\Mux24~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~13 .lut_mask = 16'hF388;
defparam \Mux24~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N1
dffeas \regs[3][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][7] .is_wysiwyg = "true";
defparam \regs[3][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N0
cycloneive_lcell_comb \Mux24~14 (
// Equation(s):
// \Mux24~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][7]~q ))) # (!dcifimemload_22 & (\regs[1][7]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[1][7]~q ),
	.datac(\regs[3][7]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux24~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~14 .lut_mask = 16'hA088;
defparam \Mux24~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N16
cycloneive_lcell_comb \Mux24~15 (
// Equation(s):
// \Mux24~15_combout  = (\Mux24~14_combout ) # ((dcifimemload_22 & (\regs[2][7]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\regs[2][7]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux24~14_combout ),
	.cin(gnd),
	.combout(\Mux24~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~15 .lut_mask = 16'hFF08;
defparam \Mux24~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N10
cycloneive_lcell_comb \Mux24~16 (
// Equation(s):
// \Mux24~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & (\Mux24~13_combout )) # (!dcifimemload_23 & ((\Mux24~15_combout )))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux24~13_combout ),
	.datad(\Mux24~15_combout ),
	.cin(gnd),
	.combout(\Mux24~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~16 .lut_mask = 16'hD9C8;
defparam \Mux24~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N20
cycloneive_lcell_comb \Mux24~19 (
// Equation(s):
// \Mux24~19_combout  = (dcifimemload_24 & ((\Mux24~16_combout  & ((\Mux24~18_combout ))) # (!\Mux24~16_combout  & (\Mux24~11_combout )))) # (!dcifimemload_24 & (((\Mux24~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux24~11_combout ),
	.datac(\Mux24~18_combout ),
	.datad(\Mux24~16_combout ),
	.cin(gnd),
	.combout(\Mux24~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~19 .lut_mask = 16'hF588;
defparam \Mux24~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N10
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[21][7]~q )) # (!dcifimemload_23 & ((\regs[17][7]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[21][7]~q ),
	.datac(\regs[17][7]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hEE50;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N20
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (dcifimemload_24 & ((\Mux24~0_combout  & ((\regs[29][7]~q ))) # (!\Mux24~0_combout  & (\regs[25][7]~q )))) # (!dcifimemload_24 & (((\Mux24~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[25][7]~q ),
	.datac(\regs[29][7]~q ),
	.datad(\Mux24~0_combout ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hF588;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y44_N25
dffeas \regs[28][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][7] .is_wysiwyg = "true";
defparam \regs[28][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N21
dffeas \regs[16][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][7] .is_wysiwyg = "true";
defparam \regs[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N30
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (dcifimemload_24 & ((\regs[24][7]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[16][7]~q  & !dcifimemload_23))))

	.dataa(\regs[24][7]~q ),
	.datab(\regs[16][7]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hF0AC;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N12
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (\Mux24~4_combout  & (((\regs[28][7]~q ) # (!dcifimemload_23)))) # (!\Mux24~4_combout  & (\regs[20][7]~q  & ((dcifimemload_23))))

	.dataa(\regs[20][7]~q ),
	.datab(\regs[28][7]~q ),
	.datac(\Mux24~4_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hCAF0;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N31
dffeas \regs[22][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~49_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][7] .is_wysiwyg = "true";
defparam \regs[22][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N16
cycloneive_lcell_comb \regs[18][7]~feeder (
// Equation(s):
// \regs[18][7]~feeder_combout  = \regs~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~49_combout ),
	.cin(gnd),
	.combout(\regs[18][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[18][7]~feeder .lut_mask = 16'hFF00;
defparam \regs[18][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N17
dffeas \regs[18][7] (
	.clk(CLK),
	.d(\regs[18][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][7] .is_wysiwyg = "true";
defparam \regs[18][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N14
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (dcifimemload_24 & ((\regs[26][7]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[18][7]~q  & !dcifimemload_23))))

	.dataa(\regs[26][7]~q ),
	.datab(\regs[18][7]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'hF0AC;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N30
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (\Mux24~2_combout  & ((\regs[30][7]~q ) # ((!dcifimemload_23)))) # (!\Mux24~2_combout  & (((\regs[22][7]~q  & dcifimemload_23))))

	.dataa(\regs[30][7]~q ),
	.datab(\regs[22][7]~q ),
	.datac(\Mux24~2_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'hACF0;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N4
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux24~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux24~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux24~5_combout ),
	.datad(\Mux24~3_combout ),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hBA98;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N16
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[23][7]~q )) # (!dcifimemload_23 & ((\regs[19][7]~q )))))

	.dataa(\regs[23][7]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[19][7]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'hEE30;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N30
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (dcifimemload_24 & ((\Mux24~7_combout  & ((\regs[31][7]~q ))) # (!\Mux24~7_combout  & (\regs[27][7]~q )))) # (!dcifimemload_24 & (((\Mux24~7_combout ))))

	.dataa(\regs[27][7]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[31][7]~q ),
	.datad(\Mux24~7_combout ),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'hF388;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y45_N6
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// \Mux24~9_combout  = (dcifimemload_21 & ((\Mux24~6_combout  & ((\Mux24~8_combout ))) # (!\Mux24~6_combout  & (\Mux24~1_combout )))) # (!dcifimemload_21 & (((\Mux24~6_combout ))))

	.dataa(\Mux24~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux24~6_combout ),
	.datad(\Mux24~8_combout ),
	.cin(gnd),
	.combout(\Mux24~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hF838;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N28
cycloneive_lcell_comb \regs~50 (
// Equation(s):
// \regs~50_combout  = (\Add1~8_combout  & (!cuifRegSel_0 & cuifRegSel_11))

	.dataa(Add14),
	.datab(cuifRegSel_0),
	.datac(gnd),
	.datad(cuifRegSel_11),
	.cin(gnd),
	.combout(\regs~50_combout ),
	.cout());
// synopsys translate_off
defparam \regs~50 .lut_mask = 16'h2200;
defparam \regs~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N16
cycloneive_lcell_comb \regs~51 (
// Equation(s):
// \regs~51_combout  = (cuifRegSel_0 & (((ramiframload_6)))) # (!cuifRegSel_0 & (!Selector0 & ((Mux251))))

	.dataa(Selector0),
	.datab(ramiframload_6),
	.datac(cuifRegSel_0),
	.datad(Mux251),
	.cin(gnd),
	.combout(\regs~51_combout ),
	.cout());
// synopsys translate_off
defparam \regs~51 .lut_mask = 16'hC5C0;
defparam \regs~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N12
cycloneive_lcell_comb \regs~52 (
// Equation(s):
// \regs~52_combout  = (!\Equal0~1_combout  & ((\regs~50_combout ) # ((!cuifRegSel_11 & \regs~51_combout ))))

	.dataa(\Equal0~1_combout ),
	.datab(cuifRegSel_11),
	.datac(\regs~50_combout ),
	.datad(\regs~51_combout ),
	.cin(gnd),
	.combout(\regs~52_combout ),
	.cout());
// synopsys translate_off
defparam \regs~52 .lut_mask = 16'h5150;
defparam \regs~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N13
dffeas \regs[25][6] (
	.clk(CLK),
	.d(\regs~52_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][6] .is_wysiwyg = "true";
defparam \regs[25][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N26
cycloneive_lcell_comb \regs[29][6]~feeder (
// Equation(s):
// \regs[29][6]~feeder_combout  = \regs~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[29][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[29][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N27
dffeas \regs[29][6] (
	.clk(CLK),
	.d(\regs[29][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][6] .is_wysiwyg = "true";
defparam \regs[29][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N9
dffeas \regs[21][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][6] .is_wysiwyg = "true";
defparam \regs[21][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N8
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (dcifimemload_18 & (((\regs[21][6]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[17][6]~q  & ((!dcifimemload_19))))

	.dataa(\regs[17][6]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[21][6]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hCCE2;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N10
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (\Mux57~0_combout  & (((\regs[29][6]~q ) # (!dcifimemload_19)))) # (!\Mux57~0_combout  & (\regs[25][6]~q  & ((dcifimemload_19))))

	.dataa(\regs[25][6]~q ),
	.datab(\regs[29][6]~q ),
	.datac(\Mux57~0_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hCAF0;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N5
dffeas \regs[31][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][6] .is_wysiwyg = "true";
defparam \regs[31][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N4
cycloneive_lcell_comb \regs[27][6]~feeder (
// Equation(s):
// \regs[27][6]~feeder_combout  = \regs~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~52_combout ),
	.cin(gnd),
	.combout(\regs[27][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][6]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N5
dffeas \regs[27][6] (
	.clk(CLK),
	.d(\regs[27][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][6] .is_wysiwyg = "true";
defparam \regs[27][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N16
cycloneive_lcell_comb \regs[23][6]~feeder (
// Equation(s):
// \regs[23][6]~feeder_combout  = \regs~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[23][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[23][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N17
dffeas \regs[23][6] (
	.clk(CLK),
	.d(\regs[23][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][6] .is_wysiwyg = "true";
defparam \regs[23][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N6
cycloneive_lcell_comb \Mux57~7 (
// Equation(s):
// \Mux57~7_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\regs[23][6]~q ))) # (!dcifimemload_18 & (\regs[19][6]~q ))))

	.dataa(\regs[19][6]~q ),
	.datab(\regs[23][6]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux57~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~7 .lut_mask = 16'hFC0A;
defparam \Mux57~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N0
cycloneive_lcell_comb \Mux57~8 (
// Equation(s):
// \Mux57~8_combout  = (dcifimemload_19 & ((\Mux57~7_combout  & (\regs[31][6]~q )) # (!\Mux57~7_combout  & ((\regs[27][6]~q ))))) # (!dcifimemload_19 & (((\Mux57~7_combout ))))

	.dataa(\regs[31][6]~q ),
	.datab(\regs[27][6]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux57~7_combout ),
	.cin(gnd),
	.combout(\Mux57~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~8 .lut_mask = 16'hAFC0;
defparam \Mux57~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N29
dffeas \regs[22][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][6] .is_wysiwyg = "true";
defparam \regs[22][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N17
dffeas \regs[30][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][6] .is_wysiwyg = "true";
defparam \regs[30][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N28
cycloneive_lcell_comb \Mux57~3 (
// Equation(s):
// \Mux57~3_combout  = (\Mux57~2_combout  & (((\regs[30][6]~q )) # (!dcifimemload_18))) # (!\Mux57~2_combout  & (dcifimemload_18 & (\regs[22][6]~q )))

	.dataa(\Mux57~2_combout ),
	.datab(dcifimemload_18),
	.datac(\regs[22][6]~q ),
	.datad(\regs[30][6]~q ),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~3 .lut_mask = 16'hEA62;
defparam \Mux57~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N25
dffeas \regs[28][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][6] .is_wysiwyg = "true";
defparam \regs[28][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N13
dffeas \regs[20][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][6] .is_wysiwyg = "true";
defparam \regs[20][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N19
dffeas \regs[16][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][6] .is_wysiwyg = "true";
defparam \regs[16][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N7
dffeas \regs[24][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][6] .is_wysiwyg = "true";
defparam \regs[24][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N6
cycloneive_lcell_comb \Mux57~4 (
// Equation(s):
// \Mux57~4_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[24][6]~q ))) # (!dcifimemload_19 & (\regs[16][6]~q ))))

	.dataa(dcifimemload_18),
	.datab(\regs[16][6]~q ),
	.datac(\regs[24][6]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~4 .lut_mask = 16'hFA44;
defparam \Mux57~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N12
cycloneive_lcell_comb \Mux57~5 (
// Equation(s):
// \Mux57~5_combout  = (dcifimemload_18 & ((\Mux57~4_combout  & (\regs[28][6]~q )) # (!\Mux57~4_combout  & ((\regs[20][6]~q ))))) # (!dcifimemload_18 & (((\Mux57~4_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[28][6]~q ),
	.datac(\regs[20][6]~q ),
	.datad(\Mux57~4_combout ),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~5 .lut_mask = 16'hDDA0;
defparam \Mux57~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N20
cycloneive_lcell_comb \Mux57~6 (
// Equation(s):
// \Mux57~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux57~3_combout )) # (!dcifimemload_17 & ((\Mux57~5_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux57~3_combout ),
	.datad(\Mux57~5_combout ),
	.cin(gnd),
	.combout(\Mux57~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~6 .lut_mask = 16'hD9C8;
defparam \Mux57~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N25
dffeas \regs[14][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][6] .is_wysiwyg = "true";
defparam \regs[14][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N31
dffeas \regs[15][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][6] .is_wysiwyg = "true";
defparam \regs[15][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N9
dffeas \regs[13][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][6] .is_wysiwyg = "true";
defparam \regs[13][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N11
dffeas \regs[12][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][6] .is_wysiwyg = "true";
defparam \regs[12][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N10
cycloneive_lcell_comb \Mux57~17 (
// Equation(s):
// \Mux57~17_combout  = (dcifimemload_16 & ((\regs[13][6]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[12][6]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[13][6]~q ),
	.datac(\regs[12][6]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux57~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~17 .lut_mask = 16'hAAD8;
defparam \Mux57~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N30
cycloneive_lcell_comb \Mux57~18 (
// Equation(s):
// \Mux57~18_combout  = (dcifimemload_17 & ((\Mux57~17_combout  & ((\regs[15][6]~q ))) # (!\Mux57~17_combout  & (\regs[14][6]~q )))) # (!dcifimemload_17 & (((\Mux57~17_combout ))))

	.dataa(\regs[14][6]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[15][6]~q ),
	.datad(\Mux57~17_combout ),
	.cin(gnd),
	.combout(\Mux57~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~18 .lut_mask = 16'hF388;
defparam \Mux57~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N17
dffeas \regs[11][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][6] .is_wysiwyg = "true";
defparam \regs[11][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N29
dffeas \regs[9][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][6] .is_wysiwyg = "true";
defparam \regs[9][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N7
dffeas \regs[10][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][6] .is_wysiwyg = "true";
defparam \regs[10][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N6
cycloneive_lcell_comb \Mux57~10 (
// Equation(s):
// \Mux57~10_combout  = (dcifimemload_17 & (((\regs[10][6]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\regs[8][6]~q  & ((!dcifimemload_16))))

	.dataa(\regs[8][6]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[10][6]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux57~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~10 .lut_mask = 16'hCCE2;
defparam \Mux57~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N28
cycloneive_lcell_comb \Mux57~11 (
// Equation(s):
// \Mux57~11_combout  = (dcifimemload_16 & ((\Mux57~10_combout  & (\regs[11][6]~q )) # (!\Mux57~10_combout  & ((\regs[9][6]~q ))))) # (!dcifimemload_16 & (((\Mux57~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[11][6]~q ),
	.datac(\regs[9][6]~q ),
	.datad(\Mux57~10_combout ),
	.cin(gnd),
	.combout(\Mux57~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~11 .lut_mask = 16'hDDA0;
defparam \Mux57~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y32_N11
dffeas \regs[2][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][6] .is_wysiwyg = "true";
defparam \regs[2][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N27
dffeas \regs[3][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][6] .is_wysiwyg = "true";
defparam \regs[3][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N25
dffeas \regs[1][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][6] .is_wysiwyg = "true";
defparam \regs[1][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N24
cycloneive_lcell_comb \Mux57~14 (
// Equation(s):
// \Mux57~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][6]~q )) # (!dcifimemload_17 & ((\regs[1][6]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[3][6]~q ),
	.datac(\regs[1][6]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux57~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~14 .lut_mask = 16'h88A0;
defparam \Mux57~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N10
cycloneive_lcell_comb \Mux57~15 (
// Equation(s):
// \Mux57~15_combout  = (\Mux57~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][6]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][6]~q ),
	.datad(\Mux57~14_combout ),
	.cin(gnd),
	.combout(\Mux57~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~15 .lut_mask = 16'hFF40;
defparam \Mux57~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N18
cycloneive_lcell_comb \regs[6][6]~feeder (
// Equation(s):
// \regs[6][6]~feeder_combout  = \regs~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[6][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[6][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N19
dffeas \regs[6][6] (
	.clk(CLK),
	.d(\regs[6][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][6] .is_wysiwyg = "true";
defparam \regs[6][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N23
dffeas \regs[7][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][6] .is_wysiwyg = "true";
defparam \regs[7][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N3
dffeas \regs[4][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][6] .is_wysiwyg = "true";
defparam \regs[4][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N16
cycloneive_lcell_comb \Mux57~12 (
// Equation(s):
// \Mux57~12_combout  = (dcifimemload_16 & ((\regs[5][6]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][6]~q  & !dcifimemload_17))))

	.dataa(\regs[5][6]~q ),
	.datab(\regs[4][6]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux57~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~12 .lut_mask = 16'hF0AC;
defparam \Mux57~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N22
cycloneive_lcell_comb \Mux57~13 (
// Equation(s):
// \Mux57~13_combout  = (dcifimemload_17 & ((\Mux57~12_combout  & ((\regs[7][6]~q ))) # (!\Mux57~12_combout  & (\regs[6][6]~q )))) # (!dcifimemload_17 & (((\Mux57~12_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][6]~q ),
	.datac(\regs[7][6]~q ),
	.datad(\Mux57~12_combout ),
	.cin(gnd),
	.combout(\Mux57~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~13 .lut_mask = 16'hF588;
defparam \Mux57~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N28
cycloneive_lcell_comb \Mux57~16 (
// Equation(s):
// \Mux57~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux57~13_combout ))) # (!dcifimemload_18 & (\Mux57~15_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux57~15_combout ),
	.datad(\Mux57~13_combout ),
	.cin(gnd),
	.combout(\Mux57~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~16 .lut_mask = 16'hDC98;
defparam \Mux57~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N19
dffeas \regs[19][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][6] .is_wysiwyg = "true";
defparam \regs[19][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N18
cycloneive_lcell_comb \Mux25~7 (
// Equation(s):
// \Mux25~7_combout  = (dcifimemload_24 & ((\regs[27][6]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[19][6]~q  & !dcifimemload_23))))

	.dataa(\regs[27][6]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[19][6]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~7 .lut_mask = 16'hCCB8;
defparam \Mux25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N4
cycloneive_lcell_comb \Mux25~8 (
// Equation(s):
// \Mux25~8_combout  = (dcifimemload_23 & ((\Mux25~7_combout  & ((\regs[31][6]~q ))) # (!\Mux25~7_combout  & (\regs[23][6]~q )))) # (!dcifimemload_23 & (((\Mux25~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[23][6]~q ),
	.datac(\regs[31][6]~q ),
	.datad(\Mux25~7_combout ),
	.cin(gnd),
	.combout(\Mux25~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~8 .lut_mask = 16'hF588;
defparam \Mux25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N9
dffeas \regs[18][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][6] .is_wysiwyg = "true";
defparam \regs[18][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N8
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[22][6]~q )) # (!dcifimemload_23 & ((\regs[18][6]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[22][6]~q ),
	.datac(\regs[18][6]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'hEE50;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N16
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (\Mux25~2_combout  & (((\regs[30][6]~q ) # (!dcifimemload_24)))) # (!\Mux25~2_combout  & (\regs[26][6]~q  & ((dcifimemload_24))))

	.dataa(\regs[26][6]~q ),
	.datab(\regs[30][6]~q ),
	.datac(\Mux25~2_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hCAF0;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N30
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (dcifimemload_23 & (((\regs[20][6]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[16][6]~q  & ((!dcifimemload_24))))

	.dataa(\regs[16][6]~q ),
	.datab(\regs[20][6]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hF0CA;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N20
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (\Mux25~4_combout  & ((\regs[28][6]~q ) # ((!dcifimemload_24)))) # (!\Mux25~4_combout  & (((\regs[24][6]~q  & dcifimemload_24))))

	.dataa(\regs[28][6]~q ),
	.datab(\regs[24][6]~q ),
	.datac(\Mux25~4_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hACF0;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N8
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// \Mux25~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux25~3_combout )) # (!dcifimemload_22 & ((\Mux25~5_combout )))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux25~3_combout ),
	.datad(\Mux25~5_combout ),
	.cin(gnd),
	.combout(\Mux25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hD9C8;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N8
cycloneive_lcell_comb \regs[17][6]~feeder (
// Equation(s):
// \regs[17][6]~feeder_combout  = \regs~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~52_combout ),
	.cin(gnd),
	.combout(\regs[17][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][6]~feeder .lut_mask = 16'hFF00;
defparam \regs[17][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N9
dffeas \regs[17][6] (
	.clk(CLK),
	.d(\regs[17][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][6] .is_wysiwyg = "true";
defparam \regs[17][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N22
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (dcifimemload_24 & ((\regs[25][6]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[17][6]~q  & !dcifimemload_23))))

	.dataa(\regs[25][6]~q ),
	.datab(\regs[17][6]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hF0AC;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N20
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Mux25~0_combout  & (((\regs[29][6]~q ) # (!dcifimemload_23)))) # (!\Mux25~0_combout  & (\regs[21][6]~q  & ((dcifimemload_23))))

	.dataa(\regs[21][6]~q ),
	.datab(\regs[29][6]~q ),
	.datac(\Mux25~0_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hCAF0;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N22
cycloneive_lcell_comb \Mux25~9 (
// Equation(s):
// \Mux25~9_combout  = (dcifimemload_21 & ((\Mux25~6_combout  & (\Mux25~8_combout )) # (!\Mux25~6_combout  & ((\Mux25~1_combout ))))) # (!dcifimemload_21 & (((\Mux25~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux25~8_combout ),
	.datac(\Mux25~6_combout ),
	.datad(\Mux25~1_combout ),
	.cin(gnd),
	.combout(\Mux25~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~9 .lut_mask = 16'hDAD0;
defparam \Mux25~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N29
dffeas \regs[5][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][6] .is_wysiwyg = "true";
defparam \regs[5][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \Mux25~10 (
// Equation(s):
// \Mux25~10_combout  = (dcifimemload_21 & (((\regs[5][6]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][6]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][6]~q ),
	.datac(\regs[5][6]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux25~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~10 .lut_mask = 16'hAAE4;
defparam \Mux25~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N12
cycloneive_lcell_comb \Mux25~11 (
// Equation(s):
// \Mux25~11_combout  = (dcifimemload_22 & ((\Mux25~10_combout  & ((\regs[7][6]~q ))) # (!\Mux25~10_combout  & (\regs[6][6]~q )))) # (!dcifimemload_22 & (((\Mux25~10_combout ))))

	.dataa(\regs[6][6]~q ),
	.datab(\regs[7][6]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux25~10_combout ),
	.cin(gnd),
	.combout(\Mux25~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~11 .lut_mask = 16'hCFA0;
defparam \Mux25~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N8
cycloneive_lcell_comb \Mux25~17 (
// Equation(s):
// \Mux25~17_combout  = (dcifimemload_21 & (((\regs[13][6]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][6]~q  & ((!dcifimemload_22))))

	.dataa(\regs[12][6]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[13][6]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux25~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~17 .lut_mask = 16'hCCE2;
defparam \Mux25~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N24
cycloneive_lcell_comb \Mux25~18 (
// Equation(s):
// \Mux25~18_combout  = (dcifimemload_22 & ((\Mux25~17_combout  & (\regs[15][6]~q )) # (!\Mux25~17_combout  & ((\regs[14][6]~q ))))) # (!dcifimemload_22 & (((\Mux25~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][6]~q ),
	.datac(\regs[14][6]~q ),
	.datad(\Mux25~17_combout ),
	.cin(gnd),
	.combout(\Mux25~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~18 .lut_mask = 16'hDDA0;
defparam \Mux25~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N26
cycloneive_lcell_comb \Mux25~14 (
// Equation(s):
// \Mux25~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][6]~q ))) # (!dcifimemload_22 & (\regs[1][6]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[1][6]~q ),
	.datac(\regs[3][6]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux25~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~14 .lut_mask = 16'hA088;
defparam \Mux25~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N4
cycloneive_lcell_comb \Mux25~15 (
// Equation(s):
// \Mux25~15_combout  = (\Mux25~14_combout ) # ((\regs[2][6]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\regs[2][6]~q ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux25~14_combout ),
	.cin(gnd),
	.combout(\Mux25~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~15 .lut_mask = 16'hFF08;
defparam \Mux25~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N18
cycloneive_lcell_comb \Mux25~12 (
// Equation(s):
// \Mux25~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][6]~q ))) # (!dcifimemload_22 & (\regs[8][6]~q ))))

	.dataa(\regs[8][6]~q ),
	.datab(\regs[10][6]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux25~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~12 .lut_mask = 16'hFC0A;
defparam \Mux25~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N16
cycloneive_lcell_comb \Mux25~13 (
// Equation(s):
// \Mux25~13_combout  = (dcifimemload_21 & ((\Mux25~12_combout  & ((\regs[11][6]~q ))) # (!\Mux25~12_combout  & (\regs[9][6]~q )))) # (!dcifimemload_21 & (((\Mux25~12_combout ))))

	.dataa(\regs[9][6]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[11][6]~q ),
	.datad(\Mux25~12_combout ),
	.cin(gnd),
	.combout(\Mux25~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~13 .lut_mask = 16'hF388;
defparam \Mux25~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N6
cycloneive_lcell_comb \Mux25~16 (
// Equation(s):
// \Mux25~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & ((\Mux25~13_combout ))) # (!dcifimemload_24 & (\Mux25~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux25~15_combout ),
	.datad(\Mux25~13_combout ),
	.cin(gnd),
	.combout(\Mux25~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~16 .lut_mask = 16'hDC98;
defparam \Mux25~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N20
cycloneive_lcell_comb \Mux25~19 (
// Equation(s):
// \Mux25~19_combout  = (dcifimemload_23 & ((\Mux25~16_combout  & ((\Mux25~18_combout ))) # (!\Mux25~16_combout  & (\Mux25~11_combout )))) # (!dcifimemload_23 & (((\Mux25~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux25~11_combout ),
	.datac(\Mux25~18_combout ),
	.datad(\Mux25~16_combout ),
	.cin(gnd),
	.combout(\Mux25~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~19 .lut_mask = 16'hF588;
defparam \Mux25~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N14
cycloneive_lcell_comb \regs~53 (
// Equation(s):
// \regs~53_combout  = (!cuifRegSel_0 & (\Add1~6_combout  & cuifRegSel_11))

	.dataa(cuifRegSel_0),
	.datab(Add13),
	.datac(gnd),
	.datad(cuifRegSel_11),
	.cin(gnd),
	.combout(\regs~53_combout ),
	.cout());
// synopsys translate_off
defparam \regs~53 .lut_mask = 16'h4400;
defparam \regs~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N6
cycloneive_lcell_comb \regs~54 (
// Equation(s):
// \regs~54_combout  = (cuifRegSel_0 & (ramiframload_51)) # (!cuifRegSel_0 & (((Mux261 & !Selector0))))

	.dataa(ramiframload_5),
	.datab(cuifRegSel_0),
	.datac(Mux261),
	.datad(Selector0),
	.cin(gnd),
	.combout(\regs~54_combout ),
	.cout());
// synopsys translate_off
defparam \regs~54 .lut_mask = 16'h88B8;
defparam \regs~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N26
cycloneive_lcell_comb \regs~55 (
// Equation(s):
// \regs~55_combout  = (!\Equal0~1_combout  & ((\regs~53_combout ) # ((!cuifRegSel_11 & \regs~54_combout ))))

	.dataa(\Equal0~1_combout ),
	.datab(cuifRegSel_11),
	.datac(\regs~53_combout ),
	.datad(\regs~54_combout ),
	.cin(gnd),
	.combout(\regs~55_combout ),
	.cout());
// synopsys translate_off
defparam \regs~55 .lut_mask = 16'h5150;
defparam \regs~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N6
cycloneive_lcell_comb \regs[23][5]~feeder (
// Equation(s):
// \regs[23][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[23][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N7
dffeas \regs[23][5] (
	.clk(CLK),
	.d(\regs[23][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][5] .is_wysiwyg = "true";
defparam \regs[23][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N28
cycloneive_lcell_comb \regs[27][5]~feeder (
// Equation(s):
// \regs[27][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[27][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N29
dffeas \regs[27][5] (
	.clk(CLK),
	.d(\regs[27][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][5] .is_wysiwyg = "true";
defparam \regs[27][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N30
cycloneive_lcell_comb \Mux58~7 (
// Equation(s):
// \Mux58~7_combout  = (dcifimemload_19 & (((\regs[27][5]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\regs[19][5]~q  & ((!dcifimemload_18))))

	.dataa(\regs[19][5]~q ),
	.datab(\regs[27][5]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux58~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~7 .lut_mask = 16'hF0CA;
defparam \Mux58~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N9
dffeas \regs[31][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][5] .is_wysiwyg = "true";
defparam \regs[31][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N16
cycloneive_lcell_comb \Mux58~8 (
// Equation(s):
// \Mux58~8_combout  = (dcifimemload_18 & ((\Mux58~7_combout  & ((\regs[31][5]~q ))) # (!\Mux58~7_combout  & (\regs[23][5]~q )))) # (!dcifimemload_18 & (((\Mux58~7_combout ))))

	.dataa(\regs[23][5]~q ),
	.datab(dcifimemload_18),
	.datac(\Mux58~7_combout ),
	.datad(\regs[31][5]~q ),
	.cin(gnd),
	.combout(\Mux58~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~8 .lut_mask = 16'hF838;
defparam \Mux58~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N20
cycloneive_lcell_comb \regs[21][5]~feeder (
// Equation(s):
// \regs[21][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~55_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[21][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][5]~feeder .lut_mask = 16'hF0F0;
defparam \regs[21][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N21
dffeas \regs[21][5] (
	.clk(CLK),
	.d(\regs[21][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][5] .is_wysiwyg = "true";
defparam \regs[21][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N4
cycloneive_lcell_comb \regs[29][5]~feeder (
// Equation(s):
// \regs[29][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[29][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[29][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N5
dffeas \regs[29][5] (
	.clk(CLK),
	.d(\regs[29][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][5] .is_wysiwyg = "true";
defparam \regs[29][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N28
cycloneive_lcell_comb \regs[25][5]~feeder (
// Equation(s):
// \regs[25][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[25][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[25][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[25][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N29
dffeas \regs[25][5] (
	.clk(CLK),
	.d(\regs[25][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][5] .is_wysiwyg = "true";
defparam \regs[25][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N14
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[25][5]~q ))) # (!dcifimemload_19 & (\regs[17][5]~q ))))

	.dataa(\regs[17][5]~q ),
	.datab(\regs[25][5]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hFC0A;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N30
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (dcifimemload_18 & ((\Mux58~0_combout  & ((\regs[29][5]~q ))) # (!\Mux58~0_combout  & (\regs[21][5]~q )))) # (!dcifimemload_18 & (((\Mux58~0_combout ))))

	.dataa(dcifimemload_18),
	.datab(\regs[21][5]~q ),
	.datac(\regs[29][5]~q ),
	.datad(\Mux58~0_combout ),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hF588;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N15
dffeas \regs[22][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][5] .is_wysiwyg = "true";
defparam \regs[22][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N14
cycloneive_lcell_comb \Mux58~2 (
// Equation(s):
// \Mux58~2_combout  = (dcifimemload_18 & (((\regs[22][5]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[18][5]~q  & ((!dcifimemload_19))))

	.dataa(\regs[18][5]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[22][5]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux58~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~2 .lut_mask = 16'hCCE2;
defparam \Mux58~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N9
dffeas \regs[26][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][5] .is_wysiwyg = "true";
defparam \regs[26][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N8
cycloneive_lcell_comb \Mux58~3 (
// Equation(s):
// \Mux58~3_combout  = (\Mux58~2_combout  & ((\regs[30][5]~q ) # ((!dcifimemload_19)))) # (!\Mux58~2_combout  & (((\regs[26][5]~q  & dcifimemload_19))))

	.dataa(\regs[30][5]~q ),
	.datab(\Mux58~2_combout ),
	.datac(\regs[26][5]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux58~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~3 .lut_mask = 16'hB8CC;
defparam \Mux58~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N24
cycloneive_lcell_comb \regs[24][5]~feeder (
// Equation(s):
// \regs[24][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[24][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[24][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N25
dffeas \regs[24][5] (
	.clk(CLK),
	.d(\regs[24][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][5] .is_wysiwyg = "true";
defparam \regs[24][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N20
cycloneive_lcell_comb \regs[20][5]~feeder (
// Equation(s):
// \regs[20][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~55_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[20][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][5]~feeder .lut_mask = 16'hF0F0;
defparam \regs[20][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N21
dffeas \regs[20][5] (
	.clk(CLK),
	.d(\regs[20][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][5] .is_wysiwyg = "true";
defparam \regs[20][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N20
cycloneive_lcell_comb \Mux58~4 (
// Equation(s):
// \Mux58~4_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\regs[20][5]~q ))) # (!dcifimemload_18 & (\regs[16][5]~q ))))

	.dataa(\regs[16][5]~q ),
	.datab(\regs[20][5]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux58~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~4 .lut_mask = 16'hFC0A;
defparam \Mux58~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N10
cycloneive_lcell_comb \Mux58~5 (
// Equation(s):
// \Mux58~5_combout  = (dcifimemload_19 & ((\Mux58~4_combout  & (\regs[28][5]~q )) # (!\Mux58~4_combout  & ((\regs[24][5]~q ))))) # (!dcifimemload_19 & (((\Mux58~4_combout ))))

	.dataa(\regs[28][5]~q ),
	.datab(\regs[24][5]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux58~4_combout ),
	.cin(gnd),
	.combout(\Mux58~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~5 .lut_mask = 16'hAFC0;
defparam \Mux58~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N28
cycloneive_lcell_comb \Mux58~6 (
// Equation(s):
// \Mux58~6_combout  = (dcifimemload_17 & ((\Mux58~3_combout ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((!dcifimemload_16 & \Mux58~5_combout ))))

	.dataa(\Mux58~3_combout ),
	.datab(dcifimemload_17),
	.datac(dcifimemload_16),
	.datad(\Mux58~5_combout ),
	.cin(gnd),
	.combout(\Mux58~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~6 .lut_mask = 16'hCBC8;
defparam \Mux58~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N21
dffeas \regs[14][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][5] .is_wysiwyg = "true";
defparam \regs[14][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N7
dffeas \regs[15][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][5] .is_wysiwyg = "true";
defparam \regs[15][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N15
dffeas \regs[12][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][5] .is_wysiwyg = "true";
defparam \regs[12][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N14
cycloneive_lcell_comb \Mux58~17 (
// Equation(s):
// \Mux58~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][5]~q )) # (!dcifimemload_16 & ((\regs[12][5]~q )))))

	.dataa(\regs[13][5]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][5]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux58~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~17 .lut_mask = 16'hEE30;
defparam \Mux58~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N6
cycloneive_lcell_comb \Mux58~18 (
// Equation(s):
// \Mux58~18_combout  = (dcifimemload_17 & ((\Mux58~17_combout  & ((\regs[15][5]~q ))) # (!\Mux58~17_combout  & (\regs[14][5]~q )))) # (!dcifimemload_17 & (((\Mux58~17_combout ))))

	.dataa(\regs[14][5]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[15][5]~q ),
	.datad(\Mux58~17_combout ),
	.cin(gnd),
	.combout(\Mux58~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~18 .lut_mask = 16'hF388;
defparam \Mux58~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N12
cycloneive_lcell_comb \regs[9][5]~feeder (
// Equation(s):
// \regs[9][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[9][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N13
dffeas \regs[9][5] (
	.clk(CLK),
	.d(\regs[9][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][5] .is_wysiwyg = "true";
defparam \regs[9][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N3
dffeas \regs[11][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][5] .is_wysiwyg = "true";
defparam \regs[11][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N27
dffeas \regs[10][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][5] .is_wysiwyg = "true";
defparam \regs[10][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N21
dffeas \regs[8][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][5] .is_wysiwyg = "true";
defparam \regs[8][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N20
cycloneive_lcell_comb \Mux58~12 (
// Equation(s):
// \Mux58~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][5]~q )) # (!dcifimemload_17 & ((\regs[8][5]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][5]~q ),
	.datac(\regs[8][5]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux58~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~12 .lut_mask = 16'hEE50;
defparam \Mux58~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N2
cycloneive_lcell_comb \Mux58~13 (
// Equation(s):
// \Mux58~13_combout  = (dcifimemload_16 & ((\Mux58~12_combout  & ((\regs[11][5]~q ))) # (!\Mux58~12_combout  & (\regs[9][5]~q )))) # (!dcifimemload_16 & (((\Mux58~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][5]~q ),
	.datac(\regs[11][5]~q ),
	.datad(\Mux58~12_combout ),
	.cin(gnd),
	.combout(\Mux58~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~13 .lut_mask = 16'hF588;
defparam \Mux58~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N16
cycloneive_lcell_comb \regs[2][5]~feeder (
// Equation(s):
// \regs[2][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~55_combout ),
	.cin(gnd),
	.combout(\regs[2][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[2][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[2][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N17
dffeas \regs[2][5] (
	.clk(CLK),
	.d(\regs[2][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][5] .is_wysiwyg = "true";
defparam \regs[2][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N27
dffeas \regs[1][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][5] .is_wysiwyg = "true";
defparam \regs[1][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N26
cycloneive_lcell_comb \Mux58~14 (
// Equation(s):
// \Mux58~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][5]~q )) # (!dcifimemload_17 & ((\regs[1][5]~q )))))

	.dataa(\regs[3][5]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][5]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux58~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~14 .lut_mask = 16'h88C0;
defparam \Mux58~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N2
cycloneive_lcell_comb \Mux58~15 (
// Equation(s):
// \Mux58~15_combout  = (\Mux58~14_combout ) # ((!dcifimemload_16 & (\regs[2][5]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\regs[2][5]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux58~14_combout ),
	.cin(gnd),
	.combout(\Mux58~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~15 .lut_mask = 16'hFF40;
defparam \Mux58~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N8
cycloneive_lcell_comb \Mux58~16 (
// Equation(s):
// \Mux58~16_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux58~13_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & ((\Mux58~15_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux58~13_combout ),
	.datad(\Mux58~15_combout ),
	.cin(gnd),
	.combout(\Mux58~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~16 .lut_mask = 16'hB9A8;
defparam \Mux58~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N3
dffeas \regs[7][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][5] .is_wysiwyg = "true";
defparam \regs[7][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N17
dffeas \regs[6][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][5] .is_wysiwyg = "true";
defparam \regs[6][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N19
dffeas \regs[5][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][5] .is_wysiwyg = "true";
defparam \regs[5][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N18
cycloneive_lcell_comb \Mux58~10 (
// Equation(s):
// \Mux58~10_combout  = (dcifimemload_16 & (((\regs[5][5]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][5]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][5]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[5][5]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux58~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~10 .lut_mask = 16'hCCE2;
defparam \Mux58~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N16
cycloneive_lcell_comb \Mux58~11 (
// Equation(s):
// \Mux58~11_combout  = (dcifimemload_17 & ((\Mux58~10_combout  & (\regs[7][5]~q )) # (!\Mux58~10_combout  & ((\regs[6][5]~q ))))) # (!dcifimemload_17 & (((\Mux58~10_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[7][5]~q ),
	.datac(\regs[6][5]~q ),
	.datad(\Mux58~10_combout ),
	.cin(gnd),
	.combout(\Mux58~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~11 .lut_mask = 16'hDDA0;
defparam \Mux58~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N26
cycloneive_lcell_comb \Mux26~10 (
// Equation(s):
// \Mux26~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][5]~q ))) # (!dcifimemload_22 & (\regs[8][5]~q ))))

	.dataa(\regs[8][5]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[10][5]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux26~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~10 .lut_mask = 16'hFC22;
defparam \Mux26~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N26
cycloneive_lcell_comb \Mux26~11 (
// Equation(s):
// \Mux26~11_combout  = (dcifimemload_21 & ((\Mux26~10_combout  & ((\regs[11][5]~q ))) # (!\Mux26~10_combout  & (\regs[9][5]~q )))) # (!dcifimemload_21 & (((\Mux26~10_combout ))))

	.dataa(\regs[9][5]~q ),
	.datab(\regs[11][5]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux26~10_combout ),
	.cin(gnd),
	.combout(\Mux26~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~11 .lut_mask = 16'hCFA0;
defparam \Mux26~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y36_N25
dffeas \regs[3][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][5] .is_wysiwyg = "true";
defparam \regs[3][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N24
cycloneive_lcell_comb \Mux26~14 (
// Equation(s):
// \Mux26~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][5]~q ))) # (!dcifimemload_22 & (\regs[1][5]~q ))))

	.dataa(\regs[1][5]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[3][5]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux26~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~14 .lut_mask = 16'hE200;
defparam \Mux26~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N22
cycloneive_lcell_comb \Mux26~15 (
// Equation(s):
// \Mux26~15_combout  = (\Mux26~14_combout ) # ((dcifimemload_22 & (\regs[2][5]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\regs[2][5]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux26~14_combout ),
	.cin(gnd),
	.combout(\Mux26~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~15 .lut_mask = 16'hFF08;
defparam \Mux26~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N13
dffeas \regs[4][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][5] .is_wysiwyg = "true";
defparam \regs[4][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N12
cycloneive_lcell_comb \Mux26~12 (
// Equation(s):
// \Mux26~12_combout  = (dcifimemload_21 & ((\regs[5][5]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\regs[4][5]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[5][5]~q ),
	.datac(\regs[4][5]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux26~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~12 .lut_mask = 16'hAAD8;
defparam \Mux26~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N2
cycloneive_lcell_comb \Mux26~13 (
// Equation(s):
// \Mux26~13_combout  = (dcifimemload_22 & ((\Mux26~12_combout  & ((\regs[7][5]~q ))) # (!\Mux26~12_combout  & (\regs[6][5]~q )))) # (!dcifimemload_22 & (((\Mux26~12_combout ))))

	.dataa(\regs[6][5]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[7][5]~q ),
	.datad(\Mux26~12_combout ),
	.cin(gnd),
	.combout(\Mux26~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~13 .lut_mask = 16'hF388;
defparam \Mux26~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N4
cycloneive_lcell_comb \Mux26~16 (
// Equation(s):
// \Mux26~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux26~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & (\Mux26~15_combout )))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux26~15_combout ),
	.datad(\Mux26~13_combout ),
	.cin(gnd),
	.combout(\Mux26~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~16 .lut_mask = 16'hBA98;
defparam \Mux26~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N29
dffeas \regs[13][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][5] .is_wysiwyg = "true";
defparam \regs[13][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N28
cycloneive_lcell_comb \Mux26~17 (
// Equation(s):
// \Mux26~17_combout  = (dcifimemload_21 & (((\regs[13][5]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][5]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[12][5]~q ),
	.datac(\regs[13][5]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux26~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~17 .lut_mask = 16'hAAE4;
defparam \Mux26~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N20
cycloneive_lcell_comb \Mux26~18 (
// Equation(s):
// \Mux26~18_combout  = (dcifimemload_22 & ((\Mux26~17_combout  & (\regs[15][5]~q )) # (!\Mux26~17_combout  & ((\regs[14][5]~q ))))) # (!dcifimemload_22 & (((\Mux26~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][5]~q ),
	.datac(\regs[14][5]~q ),
	.datad(\Mux26~17_combout ),
	.cin(gnd),
	.combout(\Mux26~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~18 .lut_mask = 16'hDDA0;
defparam \Mux26~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N26
cycloneive_lcell_comb \Mux26~19 (
// Equation(s):
// \Mux26~19_combout  = (dcifimemload_24 & ((\Mux26~16_combout  & ((\Mux26~18_combout ))) # (!\Mux26~16_combout  & (\Mux26~11_combout )))) # (!dcifimemload_24 & (((\Mux26~16_combout ))))

	.dataa(\Mux26~11_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux26~16_combout ),
	.datad(\Mux26~18_combout ),
	.cin(gnd),
	.combout(\Mux26~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~19 .lut_mask = 16'hF838;
defparam \Mux26~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N0
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (\Mux26~0_combout  & ((\regs[29][5]~q ) # ((!dcifimemload_24)))) # (!\Mux26~0_combout  & (((dcifimemload_24 & \regs[25][5]~q ))))

	.dataa(\Mux26~0_combout ),
	.datab(\regs[29][5]~q ),
	.datac(dcifimemload_24),
	.datad(\regs[25][5]~q ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hDA8A;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N8
cycloneive_lcell_comb \Mux26~8 (
// Equation(s):
// \Mux26~8_combout  = (\Mux26~7_combout  & (((\regs[31][5]~q )) # (!dcifimemload_24))) # (!\Mux26~7_combout  & (dcifimemload_24 & ((\regs[27][5]~q ))))

	.dataa(\Mux26~7_combout ),
	.datab(dcifimemload_24),
	.datac(\regs[31][5]~q ),
	.datad(\regs[27][5]~q ),
	.cin(gnd),
	.combout(\Mux26~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~8 .lut_mask = 16'hE6A2;
defparam \Mux26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N5
dffeas \regs[28][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~55_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][5] .is_wysiwyg = "true";
defparam \regs[28][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N14
cycloneive_lcell_comb \regs[16][5]~feeder (
// Equation(s):
// \regs[16][5]~feeder_combout  = \regs~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~55_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[16][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[16][5]~feeder .lut_mask = 16'hF0F0;
defparam \regs[16][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N15
dffeas \regs[16][5] (
	.clk(CLK),
	.d(\regs[16][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][5] .is_wysiwyg = "true";
defparam \regs[16][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N10
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[24][5]~q )) # (!dcifimemload_24 & ((\regs[16][5]~q )))))

	.dataa(\regs[24][5]~q ),
	.datab(\regs[16][5]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'hFA0C;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N4
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (dcifimemload_23 & ((\Mux26~4_combout  & ((\regs[28][5]~q ))) # (!\Mux26~4_combout  & (\regs[20][5]~q )))) # (!dcifimemload_23 & (((\Mux26~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[20][5]~q ),
	.datac(\regs[28][5]~q ),
	.datad(\Mux26~4_combout ),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hF588;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N24
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\regs[26][5]~q ))) # (!dcifimemload_24 & (\regs[18][5]~q ))))

	.dataa(\regs[18][5]~q ),
	.datab(\regs[26][5]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'hFC0A;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N8
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (dcifimemload_23 & ((\Mux26~2_combout  & (\regs[30][5]~q )) # (!\Mux26~2_combout  & ((\regs[22][5]~q ))))) # (!dcifimemload_23 & (((\Mux26~2_combout ))))

	.dataa(\regs[30][5]~q ),
	.datab(\regs[22][5]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux26~2_combout ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hAFC0;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N28
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// \Mux26~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux26~3_combout ))) # (!dcifimemload_22 & (\Mux26~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux26~5_combout ),
	.datad(\Mux26~3_combout ),
	.cin(gnd),
	.combout(\Mux26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hDC98;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N20
cycloneive_lcell_comb \Mux26~9 (
// Equation(s):
// \Mux26~9_combout  = (dcifimemload_21 & ((\Mux26~6_combout  & ((\Mux26~8_combout ))) # (!\Mux26~6_combout  & (\Mux26~1_combout )))) # (!dcifimemload_21 & (((\Mux26~6_combout ))))

	.dataa(\Mux26~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux26~8_combout ),
	.datad(\Mux26~6_combout ),
	.cin(gnd),
	.combout(\Mux26~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~9 .lut_mask = 16'hF388;
defparam \Mux26~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N2
cycloneive_lcell_comb \regs~56 (
// Equation(s):
// \regs~56_combout  = (\Add1~4_combout  & (!cuifRegSel_0 & cuifRegSel_11))

	.dataa(Add12),
	.datab(cuifRegSel_0),
	.datac(gnd),
	.datad(cuifRegSel_11),
	.cin(gnd),
	.combout(\regs~56_combout ),
	.cout());
// synopsys translate_off
defparam \regs~56 .lut_mask = 16'h2200;
defparam \regs~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N18
cycloneive_lcell_comb \regs~57 (
// Equation(s):
// \regs~57_combout  = (cuifRegSel_0 & (((ramiframload_41)))) # (!cuifRegSel_0 & (!Selector0 & ((Mux271))))

	.dataa(Selector0),
	.datab(ramiframload_4),
	.datac(cuifRegSel_0),
	.datad(Mux271),
	.cin(gnd),
	.combout(\regs~57_combout ),
	.cout());
// synopsys translate_off
defparam \regs~57 .lut_mask = 16'hC5C0;
defparam \regs~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N6
cycloneive_lcell_comb \regs~58 (
// Equation(s):
// \regs~58_combout  = (!\Equal0~1_combout  & ((\regs~56_combout ) # ((!cuifRegSel_11 & \regs~57_combout ))))

	.dataa(\Equal0~1_combout ),
	.datab(cuifRegSel_11),
	.datac(\regs~56_combout ),
	.datad(\regs~57_combout ),
	.cin(gnd),
	.combout(\regs~58_combout ),
	.cout());
// synopsys translate_off
defparam \regs~58 .lut_mask = 16'h5150;
defparam \regs~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N30
cycloneive_lcell_comb \regs[27][4]~feeder (
// Equation(s):
// \regs[27][4]~feeder_combout  = \regs~58_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~58_combout ),
	.cin(gnd),
	.combout(\regs[27][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][4]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N31
dffeas \regs[27][4] (
	.clk(CLK),
	.d(\regs[27][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][4] .is_wysiwyg = "true";
defparam \regs[27][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N15
dffeas \regs[31][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][4] .is_wysiwyg = "true";
defparam \regs[31][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N0
cycloneive_lcell_comb \regs[23][4]~feeder (
// Equation(s):
// \regs[23][4]~feeder_combout  = \regs~58_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~58_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[23][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][4]~feeder .lut_mask = 16'hF0F0;
defparam \regs[23][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N1
dffeas \regs[23][4] (
	.clk(CLK),
	.d(\regs[23][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][4] .is_wysiwyg = "true";
defparam \regs[23][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N29
dffeas \regs[19][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][4] .is_wysiwyg = "true";
defparam \regs[19][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N6
cycloneive_lcell_comb \Mux59~7 (
// Equation(s):
// \Mux59~7_combout  = (dcifimemload_18 & ((\regs[23][4]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[19][4]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\regs[23][4]~q ),
	.datac(\regs[19][4]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux59~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~7 .lut_mask = 16'hAAD8;
defparam \Mux59~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N4
cycloneive_lcell_comb \Mux59~8 (
// Equation(s):
// \Mux59~8_combout  = (\Mux59~7_combout  & (((\regs[31][4]~q ) # (!dcifimemload_19)))) # (!\Mux59~7_combout  & (\regs[27][4]~q  & ((dcifimemload_19))))

	.dataa(\regs[27][4]~q ),
	.datab(\regs[31][4]~q ),
	.datac(\Mux59~7_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux59~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~8 .lut_mask = 16'hCAF0;
defparam \Mux59~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N5
dffeas \regs[22][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][4] .is_wysiwyg = "true";
defparam \regs[22][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N7
dffeas \regs[26][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][4] .is_wysiwyg = "true";
defparam \regs[26][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N6
cycloneive_lcell_comb \Mux59~2 (
// Equation(s):
// \Mux59~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[26][4]~q ))) # (!dcifimemload_19 & (\regs[18][4]~q ))))

	.dataa(\regs[18][4]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[26][4]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux59~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~2 .lut_mask = 16'hFC22;
defparam \Mux59~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N4
cycloneive_lcell_comb \Mux59~3 (
// Equation(s):
// \Mux59~3_combout  = (dcifimemload_18 & ((\Mux59~2_combout  & (\regs[30][4]~q )) # (!\Mux59~2_combout  & ((\regs[22][4]~q ))))) # (!dcifimemload_18 & (((\Mux59~2_combout ))))

	.dataa(\regs[30][4]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[22][4]~q ),
	.datad(\Mux59~2_combout ),
	.cin(gnd),
	.combout(\Mux59~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~3 .lut_mask = 16'hBBC0;
defparam \Mux59~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N31
dffeas \regs[28][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][4] .is_wysiwyg = "true";
defparam \regs[28][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N1
dffeas \regs[20][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][4] .is_wysiwyg = "true";
defparam \regs[20][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N0
cycloneive_lcell_comb \Mux59~5 (
// Equation(s):
// \Mux59~5_combout  = (\Mux59~4_combout  & ((\regs[28][4]~q ) # ((!dcifimemload_18)))) # (!\Mux59~4_combout  & (((\regs[20][4]~q  & dcifimemload_18))))

	.dataa(\Mux59~4_combout ),
	.datab(\regs[28][4]~q ),
	.datac(\regs[20][4]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux59~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~5 .lut_mask = 16'hD8AA;
defparam \Mux59~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N4
cycloneive_lcell_comb \Mux59~6 (
// Equation(s):
// \Mux59~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux59~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & ((\Mux59~5_combout ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux59~3_combout ),
	.datad(\Mux59~5_combout ),
	.cin(gnd),
	.combout(\Mux59~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~6 .lut_mask = 16'hB9A8;
defparam \Mux59~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N7
dffeas \regs[25][4] (
	.clk(CLK),
	.d(\regs~58_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][4] .is_wysiwyg = "true";
defparam \regs[25][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N15
dffeas \regs[29][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][4] .is_wysiwyg = "true";
defparam \regs[29][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N27
dffeas \regs[21][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][4] .is_wysiwyg = "true";
defparam \regs[21][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N26
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (dcifimemload_18 & (((\regs[21][4]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[17][4]~q  & ((!dcifimemload_19))))

	.dataa(\regs[17][4]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[21][4]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hCCE2;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N2
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (\Mux59~0_combout  & (((\regs[29][4]~q ) # (!dcifimemload_19)))) # (!\Mux59~0_combout  & (\regs[25][4]~q  & ((dcifimemload_19))))

	.dataa(\regs[25][4]~q ),
	.datab(\regs[29][4]~q ),
	.datac(\Mux59~0_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hCAF0;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N11
dffeas \regs[15][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][4] .is_wysiwyg = "true";
defparam \regs[15][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N1
dffeas \regs[14][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][4] .is_wysiwyg = "true";
defparam \regs[14][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N3
dffeas \regs[12][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][4] .is_wysiwyg = "true";
defparam \regs[12][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N25
dffeas \regs[13][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][4] .is_wysiwyg = "true";
defparam \regs[13][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N24
cycloneive_lcell_comb \Mux59~17 (
// Equation(s):
// \Mux59~17_combout  = (dcifimemload_16 & (((\regs[13][4]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[12][4]~q  & ((!dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\regs[12][4]~q ),
	.datac(\regs[13][4]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux59~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~17 .lut_mask = 16'hAAE4;
defparam \Mux59~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N0
cycloneive_lcell_comb \Mux59~18 (
// Equation(s):
// \Mux59~18_combout  = (dcifimemload_17 & ((\Mux59~17_combout  & (\regs[15][4]~q )) # (!\Mux59~17_combout  & ((\regs[14][4]~q ))))) # (!dcifimemload_17 & (((\Mux59~17_combout ))))

	.dataa(\regs[15][4]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[14][4]~q ),
	.datad(\Mux59~17_combout ),
	.cin(gnd),
	.combout(\Mux59~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~18 .lut_mask = 16'hBBC0;
defparam \Mux59~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N23
dffeas \regs[10][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][4] .is_wysiwyg = "true";
defparam \regs[10][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N22
cycloneive_lcell_comb \Mux59~10 (
// Equation(s):
// \Mux59~10_combout  = (dcifimemload_17 & (((\regs[10][4]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\regs[8][4]~q  & ((!dcifimemload_16))))

	.dataa(\regs[8][4]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[10][4]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux59~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~10 .lut_mask = 16'hCCE2;
defparam \Mux59~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N5
dffeas \regs[11][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][4] .is_wysiwyg = "true";
defparam \regs[11][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N21
dffeas \regs[9][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][4] .is_wysiwyg = "true";
defparam \regs[9][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N20
cycloneive_lcell_comb \Mux59~11 (
// Equation(s):
// \Mux59~11_combout  = (\Mux59~10_combout  & ((\regs[11][4]~q ) # ((!dcifimemload_16)))) # (!\Mux59~10_combout  & (((\regs[9][4]~q  & dcifimemload_16))))

	.dataa(\Mux59~10_combout ),
	.datab(\regs[11][4]~q ),
	.datac(\regs[9][4]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux59~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~11 .lut_mask = 16'hD8AA;
defparam \Mux59~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N23
dffeas \regs[1][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][4] .is_wysiwyg = "true";
defparam \regs[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N1
dffeas \regs[3][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][4] .is_wysiwyg = "true";
defparam \regs[3][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N0
cycloneive_lcell_comb \Mux59~14 (
// Equation(s):
// \Mux59~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\regs[3][4]~q ))) # (!dcifimemload_17 & (\regs[1][4]~q ))))

	.dataa(dcifimemload_17),
	.datab(\regs[1][4]~q ),
	.datac(\regs[3][4]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux59~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~14 .lut_mask = 16'hE400;
defparam \Mux59~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N27
dffeas \regs[2][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][4] .is_wysiwyg = "true";
defparam \regs[2][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N14
cycloneive_lcell_comb \Mux59~15 (
// Equation(s):
// \Mux59~15_combout  = (\Mux59~14_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][4]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux59~14_combout ),
	.datad(\regs[2][4]~q ),
	.cin(gnd),
	.combout(\Mux59~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~15 .lut_mask = 16'hF2F0;
defparam \Mux59~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N23
dffeas \regs[7][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][4] .is_wysiwyg = "true";
defparam \regs[7][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N29
dffeas \regs[6][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][4] .is_wysiwyg = "true";
defparam \regs[6][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N28
cycloneive_lcell_comb \Mux59~13 (
// Equation(s):
// \Mux59~13_combout  = (\Mux59~12_combout  & ((\regs[7][4]~q ) # ((!dcifimemload_17)))) # (!\Mux59~12_combout  & (((\regs[6][4]~q  & dcifimemload_17))))

	.dataa(\Mux59~12_combout ),
	.datab(\regs[7][4]~q ),
	.datac(\regs[6][4]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux59~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~13 .lut_mask = 16'hD8AA;
defparam \Mux59~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N24
cycloneive_lcell_comb \Mux59~16 (
// Equation(s):
// \Mux59~16_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux59~13_combout ))) # (!dcifimemload_18 & (\Mux59~15_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux59~15_combout ),
	.datad(\Mux59~13_combout ),
	.cin(gnd),
	.combout(\Mux59~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~16 .lut_mask = 16'hDC98;
defparam \Mux59~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N23
dffeas \regs[30][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][4] .is_wysiwyg = "true";
defparam \regs[30][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N15
dffeas \regs[18][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][4] .is_wysiwyg = "true";
defparam \regs[18][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N14
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[22][4]~q )) # (!dcifimemload_23 & ((\regs[18][4]~q )))))

	.dataa(dcifimemload_24),
	.datab(\regs[22][4]~q ),
	.datac(\regs[18][4]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hEE50;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N22
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (dcifimemload_24 & ((\Mux27~2_combout  & ((\regs[30][4]~q ))) # (!\Mux27~2_combout  & (\regs[26][4]~q )))) # (!dcifimemload_24 & (((\Mux27~2_combout ))))

	.dataa(\regs[26][4]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[30][4]~q ),
	.datad(\Mux27~2_combout ),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hF388;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N24
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (dcifimemload_22 & (((dcifimemload_21) # (\Mux27~3_combout )))) # (!dcifimemload_22 & (\Mux27~5_combout  & (!dcifimemload_21)))

	.dataa(\Mux27~5_combout ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hCEC2;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N28
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (dcifimemload_24 & ((\regs[27][4]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[19][4]~q  & !dcifimemload_23))))

	.dataa(\regs[27][4]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[19][4]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'hCCB8;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N14
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (dcifimemload_23 & ((\Mux27~7_combout  & ((\regs[31][4]~q ))) # (!\Mux27~7_combout  & (\regs[23][4]~q )))) # (!dcifimemload_23 & (((\Mux27~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[23][4]~q ),
	.datac(\regs[31][4]~q ),
	.datad(\Mux27~7_combout ),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'hF588;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N25
dffeas \regs[17][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][4] .is_wysiwyg = "true";
defparam \regs[17][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N24
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (dcifimemload_24 & ((\regs[25][4]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[17][4]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[25][4]~q ),
	.datac(\regs[17][4]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hAAD8;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N14
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (dcifimemload_23 & ((\Mux27~0_combout  & ((\regs[29][4]~q ))) # (!\Mux27~0_combout  & (\regs[21][4]~q )))) # (!dcifimemload_23 & (((\Mux27~0_combout ))))

	.dataa(\regs[21][4]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[29][4]~q ),
	.datad(\Mux27~0_combout ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hF388;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N26
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// \Mux27~9_combout  = (\Mux27~6_combout  & (((\Mux27~8_combout )) # (!dcifimemload_21))) # (!\Mux27~6_combout  & (dcifimemload_21 & ((\Mux27~1_combout ))))

	.dataa(\Mux27~6_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux27~8_combout ),
	.datad(\Mux27~1_combout ),
	.cin(gnd),
	.combout(\Mux27~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hE6A2;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N2
cycloneive_lcell_comb \Mux27~17 (
// Equation(s):
// \Mux27~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\regs[13][4]~q )) # (!dcifimemload_21 & ((\regs[12][4]~q )))))

	.dataa(dcifimemload_22),
	.datab(\regs[13][4]~q ),
	.datac(\regs[12][4]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux27~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~17 .lut_mask = 16'hEE50;
defparam \Mux27~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N10
cycloneive_lcell_comb \Mux27~18 (
// Equation(s):
// \Mux27~18_combout  = (dcifimemload_22 & ((\Mux27~17_combout  & ((\regs[15][4]~q ))) # (!\Mux27~17_combout  & (\regs[14][4]~q )))) # (!dcifimemload_22 & (((\Mux27~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[14][4]~q ),
	.datac(\regs[15][4]~q ),
	.datad(\Mux27~17_combout ),
	.cin(gnd),
	.combout(\Mux27~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~18 .lut_mask = 16'hF588;
defparam \Mux27~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N1
dffeas \regs[4][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][4] .is_wysiwyg = "true";
defparam \regs[4][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N27
dffeas \regs[5][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][4] .is_wysiwyg = "true";
defparam \regs[5][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N0
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (dcifimemload_21 & ((dcifimemload_22) # ((\regs[5][4]~q )))) # (!dcifimemload_21 & (!dcifimemload_22 & (\regs[4][4]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\regs[4][4]~q ),
	.datad(\regs[5][4]~q ),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hBA98;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N22
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// \Mux27~11_combout  = (dcifimemload_22 & ((\Mux27~10_combout  & ((\regs[7][4]~q ))) # (!\Mux27~10_combout  & (\regs[6][4]~q )))) # (!dcifimemload_22 & (((\Mux27~10_combout ))))

	.dataa(\regs[6][4]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[7][4]~q ),
	.datad(\Mux27~10_combout ),
	.cin(gnd),
	.combout(\Mux27~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hF388;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N7
dffeas \regs[8][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][4] .is_wysiwyg = "true";
defparam \regs[8][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\regs[10][4]~q )) # (!dcifimemload_22 & ((\regs[8][4]~q )))))

	.dataa(dcifimemload_21),
	.datab(\regs[10][4]~q ),
	.datac(\regs[8][4]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hEE50;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N4
cycloneive_lcell_comb \Mux27~13 (
// Equation(s):
// \Mux27~13_combout  = (dcifimemload_21 & ((\Mux27~12_combout  & ((\regs[11][4]~q ))) # (!\Mux27~12_combout  & (\regs[9][4]~q )))) # (!dcifimemload_21 & (((\Mux27~12_combout ))))

	.dataa(\regs[9][4]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[11][4]~q ),
	.datad(\Mux27~12_combout ),
	.cin(gnd),
	.combout(\Mux27~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~13 .lut_mask = 16'hF388;
defparam \Mux27~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N16
cycloneive_lcell_comb \Mux27~16 (
// Equation(s):
// \Mux27~16_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\Mux27~13_combout ))) # (!dcifimemload_24 & (\Mux27~15_combout ))))

	.dataa(\Mux27~15_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux27~13_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux27~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~16 .lut_mask = 16'hFC22;
defparam \Mux27~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N2
cycloneive_lcell_comb \Mux27~19 (
// Equation(s):
// \Mux27~19_combout  = (dcifimemload_23 & ((\Mux27~16_combout  & (\Mux27~18_combout )) # (!\Mux27~16_combout  & ((\Mux27~11_combout ))))) # (!dcifimemload_23 & (((\Mux27~16_combout ))))

	.dataa(\Mux27~18_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux27~11_combout ),
	.datad(\Mux27~16_combout ),
	.cin(gnd),
	.combout(\Mux27~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~19 .lut_mask = 16'hBBC0;
defparam \Mux27~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N28
cycloneive_lcell_comb \regs~60 (
// Equation(s):
// \regs~60_combout  = (!\Equal0~1_combout  & ((\regs~59_combout ) # ((\regs~64_combout  & \Add1~2_combout ))))

	.dataa(\regs~59_combout ),
	.datab(\regs~64_combout ),
	.datac(Add11),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\regs~60_combout ),
	.cout());
// synopsys translate_off
defparam \regs~60 .lut_mask = 16'h00EA;
defparam \regs~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N23
dffeas \regs[29][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][3] .is_wysiwyg = "true";
defparam \regs[29][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N24
cycloneive_lcell_comb \regs[17][3]~feeder (
// Equation(s):
// \regs[17][3]~feeder_combout  = \regs~60_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~60_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[17][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][3]~feeder .lut_mask = 16'hF0F0;
defparam \regs[17][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N25
dffeas \regs[17][3] (
	.clk(CLK),
	.d(\regs[17][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][3] .is_wysiwyg = "true";
defparam \regs[17][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N1
dffeas \regs[25][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][3] .is_wysiwyg = "true";
defparam \regs[25][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N0
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[25][3]~q ))) # (!dcifimemload_19 & (\regs[17][3]~q ))))

	.dataa(dcifimemload_18),
	.datab(\regs[17][3]~q ),
	.datac(\regs[25][3]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hFA44;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N21
dffeas \regs[21][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][3] .is_wysiwyg = "true";
defparam \regs[21][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N6
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (\Mux60~0_combout  & ((\regs[29][3]~q ) # ((!dcifimemload_18)))) # (!\Mux60~0_combout  & (((dcifimemload_18 & \regs[21][3]~q ))))

	.dataa(\regs[29][3]~q ),
	.datab(\Mux60~0_combout ),
	.datac(dcifimemload_18),
	.datad(\regs[21][3]~q ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hBC8C;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N27
dffeas \regs[30][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][3] .is_wysiwyg = "true";
defparam \regs[30][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N25
dffeas \regs[26][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][3] .is_wysiwyg = "true";
defparam \regs[26][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N11
dffeas \regs[22][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][3] .is_wysiwyg = "true";
defparam \regs[22][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N10
cycloneive_lcell_comb \Mux60~2 (
// Equation(s):
// \Mux60~2_combout  = (dcifimemload_18 & (((\regs[22][3]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\regs[18][3]~q  & ((!dcifimemload_19))))

	.dataa(\regs[18][3]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[22][3]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~2 .lut_mask = 16'hCCE2;
defparam \Mux60~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N24
cycloneive_lcell_comb \Mux60~3 (
// Equation(s):
// \Mux60~3_combout  = (dcifimemload_19 & ((\Mux60~2_combout  & (\regs[30][3]~q )) # (!\Mux60~2_combout  & ((\regs[26][3]~q ))))) # (!dcifimemload_19 & (((\Mux60~2_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[30][3]~q ),
	.datac(\regs[26][3]~q ),
	.datad(\Mux60~2_combout ),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~3 .lut_mask = 16'hDDA0;
defparam \Mux60~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N3
dffeas \regs[28][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][3] .is_wysiwyg = "true";
defparam \regs[28][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N1
dffeas \regs[24][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][3] .is_wysiwyg = "true";
defparam \regs[24][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N0
cycloneive_lcell_comb \Mux60~5 (
// Equation(s):
// \Mux60~5_combout  = (\Mux60~4_combout  & ((\regs[28][3]~q ) # ((!dcifimemload_19)))) # (!\Mux60~4_combout  & (((\regs[24][3]~q  & dcifimemload_19))))

	.dataa(\Mux60~4_combout ),
	.datab(\regs[28][3]~q ),
	.datac(\regs[24][3]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux60~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~5 .lut_mask = 16'hD8AA;
defparam \Mux60~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N8
cycloneive_lcell_comb \Mux60~6 (
// Equation(s):
// \Mux60~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux60~3_combout )) # (!dcifimemload_17 & ((\Mux60~5_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux60~3_combout ),
	.datad(\Mux60~5_combout ),
	.cin(gnd),
	.combout(\Mux60~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~6 .lut_mask = 16'hD9C8;
defparam \Mux60~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N14
cycloneive_lcell_comb \regs[23][3]~feeder (
// Equation(s):
// \regs[23][3]~feeder_combout  = \regs~60_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~60_combout ),
	.cin(gnd),
	.combout(\regs[23][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][3]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N15
dffeas \regs[23][3] (
	.clk(CLK),
	.d(\regs[23][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][3] .is_wysiwyg = "true";
defparam \regs[23][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N3
dffeas \regs[31][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][3] .is_wysiwyg = "true";
defparam \regs[31][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N25
dffeas \regs[19][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][3] .is_wysiwyg = "true";
defparam \regs[19][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N20
cycloneive_lcell_comb \Mux60~7 (
// Equation(s):
// \Mux60~7_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[27][3]~q )) # (!dcifimemload_19 & ((\regs[19][3]~q )))))

	.dataa(\regs[27][3]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[19][3]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux60~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~7 .lut_mask = 16'hEE30;
defparam \Mux60~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N26
cycloneive_lcell_comb \Mux60~8 (
// Equation(s):
// \Mux60~8_combout  = (dcifimemload_18 & ((\Mux60~7_combout  & ((\regs[31][3]~q ))) # (!\Mux60~7_combout  & (\regs[23][3]~q )))) # (!dcifimemload_18 & (((\Mux60~7_combout ))))

	.dataa(\regs[23][3]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[31][3]~q ),
	.datad(\Mux60~7_combout ),
	.cin(gnd),
	.combout(\Mux60~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~8 .lut_mask = 16'hF388;
defparam \Mux60~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N22
cycloneive_lcell_comb \regs[14][3]~feeder (
// Equation(s):
// \regs[14][3]~feeder_combout  = \regs~60_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~60_combout ),
	.cin(gnd),
	.combout(\regs[14][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][3]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N23
dffeas \regs[14][3] (
	.clk(CLK),
	.d(\regs[14][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][3] .is_wysiwyg = "true";
defparam \regs[14][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N21
dffeas \regs[13][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][3] .is_wysiwyg = "true";
defparam \regs[13][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N20
cycloneive_lcell_comb \Mux60~17 (
// Equation(s):
// \Mux60~17_combout  = (dcifimemload_16 & (((\regs[13][3]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[12][3]~q  & ((!dcifimemload_17))))

	.dataa(\regs[12][3]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[13][3]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux60~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~17 .lut_mask = 16'hCCE2;
defparam \Mux60~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N29
dffeas \regs[15][3] (
	.clk(CLK),
	.d(\regs~60_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][3] .is_wysiwyg = "true";
defparam \regs[15][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N0
cycloneive_lcell_comb \Mux60~18 (
// Equation(s):
// \Mux60~18_combout  = (dcifimemload_17 & ((\Mux60~17_combout  & ((\regs[15][3]~q ))) # (!\Mux60~17_combout  & (\regs[14][3]~q )))) # (!dcifimemload_17 & (((\Mux60~17_combout ))))

	.dataa(\regs[14][3]~q ),
	.datab(dcifimemload_17),
	.datac(\Mux60~17_combout ),
	.datad(\regs[15][3]~q ),
	.cin(gnd),
	.combout(\Mux60~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~18 .lut_mask = 16'hF838;
defparam \Mux60~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N19
dffeas \regs[7][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][3] .is_wysiwyg = "true";
defparam \regs[7][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N1
dffeas \regs[6][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][3] .is_wysiwyg = "true";
defparam \regs[6][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N27
dffeas \regs[5][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][3] .is_wysiwyg = "true";
defparam \regs[5][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \Mux60~10 (
// Equation(s):
// \Mux60~10_combout  = (dcifimemload_16 & (((\regs[5][3]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\regs[4][3]~q  & ((!dcifimemload_17))))

	.dataa(\regs[4][3]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[5][3]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux60~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~10 .lut_mask = 16'hCCE2;
defparam \Mux60~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N0
cycloneive_lcell_comb \Mux60~11 (
// Equation(s):
// \Mux60~11_combout  = (dcifimemload_17 & ((\Mux60~10_combout  & (\regs[7][3]~q )) # (!\Mux60~10_combout  & ((\regs[6][3]~q ))))) # (!dcifimemload_17 & (((\Mux60~10_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[7][3]~q ),
	.datac(\regs[6][3]~q ),
	.datad(\Mux60~10_combout ),
	.cin(gnd),
	.combout(\Mux60~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~11 .lut_mask = 16'hDDA0;
defparam \Mux60~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N7
dffeas \regs[2][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][3] .is_wysiwyg = "true";
defparam \regs[2][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N17
dffeas \regs[3][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][3] .is_wysiwyg = "true";
defparam \regs[3][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N3
dffeas \regs[1][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][3] .is_wysiwyg = "true";
defparam \regs[1][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N16
cycloneive_lcell_comb \Mux60~14 (
// Equation(s):
// \Mux60~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][3]~q )) # (!dcifimemload_17 & ((\regs[1][3]~q )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[3][3]~q ),
	.datad(\regs[1][3]~q ),
	.cin(gnd),
	.combout(\Mux60~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~14 .lut_mask = 16'hA280;
defparam \Mux60~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N6
cycloneive_lcell_comb \Mux60~15 (
// Equation(s):
// \Mux60~15_combout  = (\Mux60~14_combout ) # ((!dcifimemload_16 & (\regs[2][3]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\regs[2][3]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux60~14_combout ),
	.cin(gnd),
	.combout(\Mux60~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~15 .lut_mask = 16'hFF40;
defparam \Mux60~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N9
dffeas \regs[11][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][3] .is_wysiwyg = "true";
defparam \regs[11][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N1
dffeas \regs[9][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][3] .is_wysiwyg = "true";
defparam \regs[9][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \regs[8][3]~feeder (
// Equation(s):
// \regs[8][3]~feeder_combout  = \regs~60_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~60_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[8][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][3]~feeder .lut_mask = 16'hF0F0;
defparam \regs[8][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N25
dffeas \regs[8][3] (
	.clk(CLK),
	.d(\regs[8][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][3] .is_wysiwyg = "true";
defparam \regs[8][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N30
cycloneive_lcell_comb \Mux60~12 (
// Equation(s):
// \Mux60~12_combout  = (dcifimemload_17 & ((\regs[10][3]~q ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((\regs[8][3]~q  & !dcifimemload_16))))

	.dataa(\regs[10][3]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[8][3]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux60~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~12 .lut_mask = 16'hCCB8;
defparam \Mux60~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N0
cycloneive_lcell_comb \Mux60~13 (
// Equation(s):
// \Mux60~13_combout  = (dcifimemload_16 & ((\Mux60~12_combout  & (\regs[11][3]~q )) # (!\Mux60~12_combout  & ((\regs[9][3]~q ))))) # (!dcifimemload_16 & (((\Mux60~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[11][3]~q ),
	.datac(\regs[9][3]~q ),
	.datad(\Mux60~12_combout ),
	.cin(gnd),
	.combout(\Mux60~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~13 .lut_mask = 16'hDDA0;
defparam \Mux60~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N20
cycloneive_lcell_comb \Mux60~16 (
// Equation(s):
// \Mux60~16_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\Mux60~13_combout ))) # (!dcifimemload_19 & (\Mux60~15_combout ))))

	.dataa(\Mux60~15_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux60~13_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux60~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~16 .lut_mask = 16'hFC22;
defparam \Mux60~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N24
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// \Mux28~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[23][3]~q )) # (!dcifimemload_23 & ((\regs[19][3]~q )))))

	.dataa(\regs[23][3]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[19][3]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hEE30;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N2
cycloneive_lcell_comb \Mux28~8 (
// Equation(s):
// \Mux28~8_combout  = (dcifimemload_24 & ((\Mux28~7_combout  & ((\regs[31][3]~q ))) # (!\Mux28~7_combout  & (\regs[27][3]~q )))) # (!dcifimemload_24 & (((\Mux28~7_combout ))))

	.dataa(\regs[27][3]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[31][3]~q ),
	.datad(\Mux28~7_combout ),
	.cin(gnd),
	.combout(\Mux28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~8 .lut_mask = 16'hF388;
defparam \Mux28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N28
cycloneive_lcell_comb \regs[18][3]~feeder (
// Equation(s):
// \regs[18][3]~feeder_combout  = \regs~60_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~60_combout ),
	.cin(gnd),
	.combout(\regs[18][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[18][3]~feeder .lut_mask = 16'hFF00;
defparam \regs[18][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N29
dffeas \regs[18][3] (
	.clk(CLK),
	.d(\regs[18][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][3] .is_wysiwyg = "true";
defparam \regs[18][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N6
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (dcifimemload_24 & ((\regs[26][3]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[18][3]~q  & !dcifimemload_23))))

	.dataa(\regs[26][3]~q ),
	.datab(\regs[18][3]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hF0AC;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N26
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (dcifimemload_23 & ((\Mux28~2_combout  & ((\regs[30][3]~q ))) # (!\Mux28~2_combout  & (\regs[22][3]~q )))) # (!dcifimemload_23 & (((\Mux28~2_combout ))))

	.dataa(\regs[22][3]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[30][3]~q ),
	.datad(\Mux28~2_combout ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hF388;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y43_N27
dffeas \regs[20][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][3] .is_wysiwyg = "true";
defparam \regs[20][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N13
dffeas \regs[16][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][3] .is_wysiwyg = "true";
defparam \regs[16][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N12
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[24][3]~q )) # (!dcifimemload_24 & ((\regs[16][3]~q )))))

	.dataa(dcifimemload_23),
	.datab(\regs[24][3]~q ),
	.datac(\regs[16][3]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hEE50;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N2
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (dcifimemload_23 & ((\Mux28~4_combout  & ((\regs[28][3]~q ))) # (!\Mux28~4_combout  & (\regs[20][3]~q )))) # (!dcifimemload_23 & (((\Mux28~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[20][3]~q ),
	.datac(\regs[28][3]~q ),
	.datad(\Mux28~4_combout ),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hF588;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N8
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux28~3_combout )) # (!dcifimemload_22 & ((\Mux28~5_combout )))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux28~3_combout ),
	.datad(\Mux28~5_combout ),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hD9C8;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N28
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (dcifimemload_23 & ((\regs[21][3]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[17][3]~q  & !dcifimemload_24))))

	.dataa(\regs[21][3]~q ),
	.datab(\regs[17][3]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hF0AC;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N22
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (dcifimemload_24 & ((\Mux28~0_combout  & ((\regs[29][3]~q ))) # (!\Mux28~0_combout  & (\regs[25][3]~q )))) # (!dcifimemload_24 & (((\Mux28~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[25][3]~q ),
	.datac(\regs[29][3]~q ),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hF588;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N14
cycloneive_lcell_comb \Mux28~9 (
// Equation(s):
// \Mux28~9_combout  = (dcifimemload_21 & ((\Mux28~6_combout  & (\Mux28~8_combout )) # (!\Mux28~6_combout  & ((\Mux28~1_combout ))))) # (!dcifimemload_21 & (((\Mux28~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux28~8_combout ),
	.datac(\Mux28~6_combout ),
	.datad(\Mux28~1_combout ),
	.cin(gnd),
	.combout(\Mux28~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~9 .lut_mask = 16'hDAD0;
defparam \Mux28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N8
cycloneive_lcell_comb \regs[10][3]~feeder (
// Equation(s):
// \regs[10][3]~feeder_combout  = \regs~60_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~60_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[10][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[10][3]~feeder .lut_mask = 16'hF0F0;
defparam \regs[10][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N9
dffeas \regs[10][3] (
	.clk(CLK),
	.d(\regs[10][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][3] .is_wysiwyg = "true";
defparam \regs[10][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N18
cycloneive_lcell_comb \Mux28~10 (
// Equation(s):
// \Mux28~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][3]~q ))) # (!dcifimemload_22 & (\regs[8][3]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][3]~q ),
	.datac(\regs[10][3]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~10 .lut_mask = 16'hFA44;
defparam \Mux28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N8
cycloneive_lcell_comb \Mux28~11 (
// Equation(s):
// \Mux28~11_combout  = (dcifimemload_21 & ((\Mux28~10_combout  & ((\regs[11][3]~q ))) # (!\Mux28~10_combout  & (\regs[9][3]~q )))) # (!dcifimemload_21 & (((\Mux28~10_combout ))))

	.dataa(\regs[9][3]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[11][3]~q ),
	.datad(\Mux28~10_combout ),
	.cin(gnd),
	.combout(\Mux28~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~11 .lut_mask = 16'hF388;
defparam \Mux28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N7
dffeas \regs[12][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][3] .is_wysiwyg = "true";
defparam \regs[12][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N6
cycloneive_lcell_comb \Mux28~17 (
// Equation(s):
// \Mux28~17_combout  = (dcifimemload_21 & ((\regs[13][3]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\regs[12][3]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[13][3]~q ),
	.datac(\regs[12][3]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux28~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~17 .lut_mask = 16'hAAD8;
defparam \Mux28~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N10
cycloneive_lcell_comb \Mux28~18 (
// Equation(s):
// \Mux28~18_combout  = (dcifimemload_22 & ((\Mux28~17_combout  & ((\regs[15][3]~q ))) # (!\Mux28~17_combout  & (\regs[14][3]~q )))) # (!dcifimemload_22 & (((\Mux28~17_combout ))))

	.dataa(\regs[14][3]~q ),
	.datab(\regs[15][3]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux28~17_combout ),
	.cin(gnd),
	.combout(\Mux28~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~18 .lut_mask = 16'hCFA0;
defparam \Mux28~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N5
dffeas \regs[4][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~60_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][3] .is_wysiwyg = "true";
defparam \regs[4][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N4
cycloneive_lcell_comb \Mux28~12 (
// Equation(s):
// \Mux28~12_combout  = (dcifimemload_21 & ((\regs[5][3]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\regs[4][3]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[5][3]~q ),
	.datac(\regs[4][3]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~12 .lut_mask = 16'hAAD8;
defparam \Mux28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N18
cycloneive_lcell_comb \Mux28~13 (
// Equation(s):
// \Mux28~13_combout  = (dcifimemload_22 & ((\Mux28~12_combout  & ((\regs[7][3]~q ))) # (!\Mux28~12_combout  & (\regs[6][3]~q )))) # (!dcifimemload_22 & (((\Mux28~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[6][3]~q ),
	.datac(\regs[7][3]~q ),
	.datad(\Mux28~12_combout ),
	.cin(gnd),
	.combout(\Mux28~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~13 .lut_mask = 16'hF588;
defparam \Mux28~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N12
cycloneive_lcell_comb \Mux28~16 (
// Equation(s):
// \Mux28~16_combout  = (dcifimemload_23 & (((dcifimemload_24) # (\Mux28~13_combout )))) # (!dcifimemload_23 & (\Mux28~15_combout  & (!dcifimemload_24)))

	.dataa(\Mux28~15_combout ),
	.datab(dcifimemload_23),
	.datac(dcifimemload_24),
	.datad(\Mux28~13_combout ),
	.cin(gnd),
	.combout(\Mux28~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~16 .lut_mask = 16'hCEC2;
defparam \Mux28~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N10
cycloneive_lcell_comb \Mux28~19 (
// Equation(s):
// \Mux28~19_combout  = (dcifimemload_24 & ((\Mux28~16_combout  & ((\Mux28~18_combout ))) # (!\Mux28~16_combout  & (\Mux28~11_combout )))) # (!dcifimemload_24 & (((\Mux28~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux28~11_combout ),
	.datac(\Mux28~18_combout ),
	.datad(\Mux28~16_combout ),
	.cin(gnd),
	.combout(\Mux28~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~19 .lut_mask = 16'hF588;
defparam \Mux28~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N4
cycloneive_lcell_comb \regs~61 (
// Equation(s):
// \regs~61_combout  = (!cuifRegSel_11 & ((cuifRegSel_0 & (ramiframload_21)) # (!cuifRegSel_0 & ((Mux291)))))

	.dataa(cuifRegSel_0),
	.datab(cuifRegSel_11),
	.datac(ramiframload_2),
	.datad(Mux291),
	.cin(gnd),
	.combout(\regs~61_combout ),
	.cout());
// synopsys translate_off
defparam \regs~61 .lut_mask = 16'h3120;
defparam \regs~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N30
cycloneive_lcell_comb \regs~62 (
// Equation(s):
// \regs~62_combout  = (!\Equal0~1_combout  & ((\regs~61_combout ) # ((\Add1~0_combout  & \regs~64_combout ))))

	.dataa(\Equal0~1_combout ),
	.datab(Add1),
	.datac(\regs~64_combout ),
	.datad(\regs~61_combout ),
	.cin(gnd),
	.combout(\regs~62_combout ),
	.cout());
// synopsys translate_off
defparam \regs~62 .lut_mask = 16'h5540;
defparam \regs~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N31
dffeas \regs[20][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][2] .is_wysiwyg = "true";
defparam \regs[20][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N1
dffeas \regs[16][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][2] .is_wysiwyg = "true";
defparam \regs[16][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N13
dffeas \regs[24][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][2] .is_wysiwyg = "true";
defparam \regs[24][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N12
cycloneive_lcell_comb \Mux61~4 (
// Equation(s):
// \Mux61~4_combout  = (dcifimemload_19 & (((\regs[24][2]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\regs[16][2]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\regs[16][2]~q ),
	.datac(\regs[24][2]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux61~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~4 .lut_mask = 16'hAAE4;
defparam \Mux61~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N30
cycloneive_lcell_comb \Mux61~5 (
// Equation(s):
// \Mux61~5_combout  = (dcifimemload_18 & ((\Mux61~4_combout  & (\regs[28][2]~q )) # (!\Mux61~4_combout  & ((\regs[20][2]~q ))))) # (!dcifimemload_18 & (((\Mux61~4_combout ))))

	.dataa(\regs[28][2]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[20][2]~q ),
	.datad(\Mux61~4_combout ),
	.cin(gnd),
	.combout(\Mux61~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~5 .lut_mask = 16'hBBC0;
defparam \Mux61~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N21
dffeas \regs[22][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][2] .is_wysiwyg = "true";
defparam \regs[22][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N19
dffeas \regs[26][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][2] .is_wysiwyg = "true";
defparam \regs[26][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N18
cycloneive_lcell_comb \Mux61~2 (
// Equation(s):
// \Mux61~2_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\regs[26][2]~q ))) # (!dcifimemload_19 & (\regs[18][2]~q ))))

	.dataa(\regs[18][2]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[26][2]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux61~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~2 .lut_mask = 16'hFC22;
defparam \Mux61~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N20
cycloneive_lcell_comb \Mux61~3 (
// Equation(s):
// \Mux61~3_combout  = (dcifimemload_18 & ((\Mux61~2_combout  & (\regs[30][2]~q )) # (!\Mux61~2_combout  & ((\regs[22][2]~q ))))) # (!dcifimemload_18 & (((\Mux61~2_combout ))))

	.dataa(\regs[30][2]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[22][2]~q ),
	.datad(\Mux61~2_combout ),
	.cin(gnd),
	.combout(\Mux61~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~3 .lut_mask = 16'hBBC0;
defparam \Mux61~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N18
cycloneive_lcell_comb \Mux61~6 (
// Equation(s):
// \Mux61~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux61~3_combout ))) # (!dcifimemload_17 & (\Mux61~5_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux61~5_combout ),
	.datad(\Mux61~3_combout ),
	.cin(gnd),
	.combout(\Mux61~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~6 .lut_mask = 16'hDC98;
defparam \Mux61~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N8
cycloneive_lcell_comb \regs[27][2]~feeder (
// Equation(s):
// \regs[27][2]~feeder_combout  = \regs~62_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~62_combout ),
	.cin(gnd),
	.combout(\regs[27][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][2]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N9
dffeas \regs[27][2] (
	.clk(CLK),
	.d(\regs[27][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][2] .is_wysiwyg = "true";
defparam \regs[27][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N28
cycloneive_lcell_comb \regs[23][2]~feeder (
// Equation(s):
// \regs[23][2]~feeder_combout  = \regs~62_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~62_combout ),
	.cin(gnd),
	.combout(\regs[23][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][2]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N29
dffeas \regs[23][2] (
	.clk(CLK),
	.d(\regs[23][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][2] .is_wysiwyg = "true";
defparam \regs[23][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N13
dffeas \regs[19][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][2] .is_wysiwyg = "true";
defparam \regs[19][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N22
cycloneive_lcell_comb \Mux61~7 (
// Equation(s):
// \Mux61~7_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[23][2]~q )) # (!dcifimemload_18 & ((\regs[19][2]~q )))))

	.dataa(dcifimemload_19),
	.datab(\regs[23][2]~q ),
	.datac(\regs[19][2]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux61~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~7 .lut_mask = 16'hEE50;
defparam \Mux61~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N11
dffeas \regs[31][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][2] .is_wysiwyg = "true";
defparam \regs[31][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N10
cycloneive_lcell_comb \Mux61~8 (
// Equation(s):
// \Mux61~8_combout  = (dcifimemload_19 & ((\Mux61~7_combout  & ((\regs[31][2]~q ))) # (!\Mux61~7_combout  & (\regs[27][2]~q )))) # (!dcifimemload_19 & (((\Mux61~7_combout ))))

	.dataa(\regs[27][2]~q ),
	.datab(dcifimemload_19),
	.datac(\Mux61~7_combout ),
	.datad(\regs[31][2]~q ),
	.cin(gnd),
	.combout(\Mux61~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~8 .lut_mask = 16'hF838;
defparam \Mux61~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N7
dffeas \regs[29][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][2] .is_wysiwyg = "true";
defparam \regs[29][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N18
cycloneive_lcell_comb \regs[25][2]~feeder (
// Equation(s):
// \regs[25][2]~feeder_combout  = \regs~62_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~62_combout ),
	.cin(gnd),
	.combout(\regs[25][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[25][2]~feeder .lut_mask = 16'hFF00;
defparam \regs[25][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N19
dffeas \regs[25][2] (
	.clk(CLK),
	.d(\regs[25][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][2] .is_wysiwyg = "true";
defparam \regs[25][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N14
cycloneive_lcell_comb \regs[17][2]~feeder (
// Equation(s):
// \regs[17][2]~feeder_combout  = \regs~62_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~62_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[17][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][2]~feeder .lut_mask = 16'hF0F0;
defparam \regs[17][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N15
dffeas \regs[17][2] (
	.clk(CLK),
	.d(\regs[17][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][2] .is_wysiwyg = "true";
defparam \regs[17][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N16
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[21][2]~q )) # (!dcifimemload_18 & ((\regs[17][2]~q )))))

	.dataa(\regs[21][2]~q ),
	.datab(\regs[17][2]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hFA0C;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N26
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (dcifimemload_19 & ((\Mux61~0_combout  & (\regs[29][2]~q )) # (!\Mux61~0_combout  & ((\regs[25][2]~q ))))) # (!dcifimemload_19 & (((\Mux61~0_combout ))))

	.dataa(\regs[29][2]~q ),
	.datab(\regs[25][2]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux61~0_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hAFC0;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N15
dffeas \regs[15][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][2] .is_wysiwyg = "true";
defparam \regs[15][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N29
dffeas \regs[14][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][2] .is_wysiwyg = "true";
defparam \regs[14][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y44_N21
dffeas \regs[13][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][2] .is_wysiwyg = "true";
defparam \regs[13][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N20
cycloneive_lcell_comb \Mux61~17 (
// Equation(s):
// \Mux61~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\regs[13][2]~q ))) # (!dcifimemload_16 & (\regs[12][2]~q ))))

	.dataa(\regs[12][2]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[13][2]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux61~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~17 .lut_mask = 16'hFC22;
defparam \Mux61~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N28
cycloneive_lcell_comb \Mux61~18 (
// Equation(s):
// \Mux61~18_combout  = (dcifimemload_17 & ((\Mux61~17_combout  & (\regs[15][2]~q )) # (!\Mux61~17_combout  & ((\regs[14][2]~q ))))) # (!dcifimemload_17 & (((\Mux61~17_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[15][2]~q ),
	.datac(\regs[14][2]~q ),
	.datad(\Mux61~17_combout ),
	.cin(gnd),
	.combout(\Mux61~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~18 .lut_mask = 16'hDDA0;
defparam \Mux61~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N19
dffeas \regs[2][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][2] .is_wysiwyg = "true";
defparam \regs[2][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N28
cycloneive_lcell_comb \regs[3][2]~feeder (
// Equation(s):
// \regs[3][2]~feeder_combout  = \regs~62_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~62_combout ),
	.cin(gnd),
	.combout(\regs[3][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][2]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N29
dffeas \regs[3][2] (
	.clk(CLK),
	.d(\regs[3][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][2] .is_wysiwyg = "true";
defparam \regs[3][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N30
cycloneive_lcell_comb \Mux61~14 (
// Equation(s):
// \Mux61~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\regs[3][2]~q ))) # (!dcifimemload_17 & (\regs[1][2]~q ))))

	.dataa(\regs[1][2]~q ),
	.datab(\regs[3][2]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux61~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~14 .lut_mask = 16'hCA00;
defparam \Mux61~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N24
cycloneive_lcell_comb \Mux61~15 (
// Equation(s):
// \Mux61~15_combout  = (\Mux61~14_combout ) # ((!dcifimemload_16 & (\regs[2][2]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\regs[2][2]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux61~14_combout ),
	.cin(gnd),
	.combout(\Mux61~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~15 .lut_mask = 16'hFF40;
defparam \Mux61~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N21
dffeas \regs[6][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][2] .is_wysiwyg = "true";
defparam \regs[6][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N11
dffeas \regs[7][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][2] .is_wysiwyg = "true";
defparam \regs[7][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N25
dffeas \regs[4][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][2] .is_wysiwyg = "true";
defparam \regs[4][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N24
cycloneive_lcell_comb \Mux61~12 (
// Equation(s):
// \Mux61~12_combout  = (dcifimemload_16 & ((\regs[5][2]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][2]~q  & !dcifimemload_17))))

	.dataa(\regs[5][2]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][2]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux61~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~12 .lut_mask = 16'hCCB8;
defparam \Mux61~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N10
cycloneive_lcell_comb \Mux61~13 (
// Equation(s):
// \Mux61~13_combout  = (dcifimemload_17 & ((\Mux61~12_combout  & ((\regs[7][2]~q ))) # (!\Mux61~12_combout  & (\regs[6][2]~q )))) # (!dcifimemload_17 & (((\Mux61~12_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[6][2]~q ),
	.datac(\regs[7][2]~q ),
	.datad(\Mux61~12_combout ),
	.cin(gnd),
	.combout(\Mux61~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~13 .lut_mask = 16'hF588;
defparam \Mux61~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N14
cycloneive_lcell_comb \Mux61~16 (
// Equation(s):
// \Mux61~16_combout  = (dcifimemload_18 & (((dcifimemload_19) # (\Mux61~13_combout )))) # (!dcifimemload_18 & (\Mux61~15_combout  & (!dcifimemload_19)))

	.dataa(dcifimemload_18),
	.datab(\Mux61~15_combout ),
	.datac(dcifimemload_19),
	.datad(\Mux61~13_combout ),
	.cin(gnd),
	.combout(\Mux61~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~16 .lut_mask = 16'hAEA4;
defparam \Mux61~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N20
cycloneive_lcell_comb \regs[9][2]~feeder (
// Equation(s):
// \regs[9][2]~feeder_combout  = \regs~62_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~62_combout ),
	.cin(gnd),
	.combout(\regs[9][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][2]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N21
dffeas \regs[9][2] (
	.clk(CLK),
	.d(\regs[9][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][2] .is_wysiwyg = "true";
defparam \regs[9][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N24
cycloneive_lcell_comb \regs[11][2]~feeder (
// Equation(s):
// \regs[11][2]~feeder_combout  = \regs~62_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~62_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[11][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][2]~feeder .lut_mask = 16'hF0F0;
defparam \regs[11][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N25
dffeas \regs[11][2] (
	.clk(CLK),
	.d(\regs[11][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][2] .is_wysiwyg = "true";
defparam \regs[11][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N22
cycloneive_lcell_comb \regs[10][2]~feeder (
// Equation(s):
// \regs[10][2]~feeder_combout  = \regs~62_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~62_combout ),
	.cin(gnd),
	.combout(\regs[10][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[10][2]~feeder .lut_mask = 16'hFF00;
defparam \regs[10][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N23
dffeas \regs[10][2] (
	.clk(CLK),
	.d(\regs[10][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][2] .is_wysiwyg = "true";
defparam \regs[10][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N24
cycloneive_lcell_comb \Mux61~10 (
// Equation(s):
// \Mux61~10_combout  = (dcifimemload_17 & (((\regs[10][2]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\regs[8][2]~q  & ((!dcifimemload_16))))

	.dataa(\regs[8][2]~q ),
	.datab(\regs[10][2]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux61~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~10 .lut_mask = 16'hF0CA;
defparam \Mux61~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N30
cycloneive_lcell_comb \Mux61~11 (
// Equation(s):
// \Mux61~11_combout  = (dcifimemload_16 & ((\Mux61~10_combout  & ((\regs[11][2]~q ))) # (!\Mux61~10_combout  & (\regs[9][2]~q )))) # (!dcifimemload_16 & (((\Mux61~10_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][2]~q ),
	.datac(\regs[11][2]~q ),
	.datad(\Mux61~10_combout ),
	.cin(gnd),
	.combout(\Mux61~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~11 .lut_mask = 16'hF588;
defparam \Mux61~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N27
dffeas \regs[28][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][2] .is_wysiwyg = "true";
defparam \regs[28][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N0
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (dcifimemload_23 & ((\regs[20][2]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[16][2]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\regs[20][2]~q ),
	.datac(\regs[16][2]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hAAD8;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N26
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (dcifimemload_24 & ((\Mux29~4_combout  & ((\regs[28][2]~q ))) # (!\Mux29~4_combout  & (\regs[24][2]~q )))) # (!dcifimemload_24 & (((\Mux29~4_combout ))))

	.dataa(\regs[24][2]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[28][2]~q ),
	.datad(\Mux29~4_combout ),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hF388;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N21
dffeas \regs[30][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][2] .is_wysiwyg = "true";
defparam \regs[30][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N17
dffeas \regs[18][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][2] .is_wysiwyg = "true";
defparam \regs[18][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N16
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[22][2]~q )) # (!dcifimemload_23 & ((\regs[18][2]~q )))))

	.dataa(\regs[22][2]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[18][2]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hEE30;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N20
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (dcifimemload_24 & ((\Mux29~2_combout  & ((\regs[30][2]~q ))) # (!\Mux29~2_combout  & (\regs[26][2]~q )))) # (!dcifimemload_24 & (((\Mux29~2_combout ))))

	.dataa(\regs[26][2]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[30][2]~q ),
	.datad(\Mux29~2_combout ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hF388;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N20
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (dcifimemload_22 & (((dcifimemload_21) # (\Mux29~3_combout )))) # (!dcifimemload_22 & (\Mux29~5_combout  & (!dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\Mux29~5_combout ),
	.datac(dcifimemload_21),
	.datad(\Mux29~3_combout ),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hAEA4;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N12
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (dcifimemload_24 & ((\regs[27][2]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\regs[19][2]~q  & !dcifimemload_23))))

	.dataa(\regs[27][2]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[19][2]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hCCB8;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N10
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (dcifimemload_23 & ((\Mux29~7_combout  & ((\regs[31][2]~q ))) # (!\Mux29~7_combout  & (\regs[23][2]~q )))) # (!dcifimemload_23 & (((\Mux29~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[23][2]~q ),
	.datac(\regs[31][2]~q ),
	.datad(\Mux29~7_combout ),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hF588;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N30
cycloneive_lcell_comb \regs[21][2]~feeder (
// Equation(s):
// \regs[21][2]~feeder_combout  = \regs~62_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~62_combout ),
	.cin(gnd),
	.combout(\regs[21][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][2]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N31
dffeas \regs[21][2] (
	.clk(CLK),
	.d(\regs[21][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][2] .is_wysiwyg = "true";
defparam \regs[21][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N30
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (dcifimemload_24 & (((\regs[25][2]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[17][2]~q  & ((!dcifimemload_23))))

	.dataa(\regs[17][2]~q ),
	.datab(dcifimemload_24),
	.datac(\regs[25][2]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hCCE2;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N6
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (dcifimemload_23 & ((\Mux29~0_combout  & ((\regs[29][2]~q ))) # (!\Mux29~0_combout  & (\regs[21][2]~q )))) # (!dcifimemload_23 & (((\Mux29~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[21][2]~q ),
	.datac(\regs[29][2]~q ),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hF588;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N30
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// \Mux29~9_combout  = (dcifimemload_21 & ((\Mux29~6_combout  & (\Mux29~8_combout )) # (!\Mux29~6_combout  & ((\Mux29~1_combout ))))) # (!dcifimemload_21 & (\Mux29~6_combout ))

	.dataa(dcifimemload_21),
	.datab(\Mux29~6_combout ),
	.datac(\Mux29~8_combout ),
	.datad(\Mux29~1_combout ),
	.cin(gnd),
	.combout(\Mux29~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hE6C4;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y44_N11
dffeas \regs[12][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][2] .is_wysiwyg = "true";
defparam \regs[12][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N10
cycloneive_lcell_comb \Mux29~17 (
// Equation(s):
// \Mux29~17_combout  = (dcifimemload_21 & ((\regs[13][2]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\regs[12][2]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[13][2]~q ),
	.datac(\regs[12][2]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux29~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~17 .lut_mask = 16'hAAD8;
defparam \Mux29~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N14
cycloneive_lcell_comb \Mux29~18 (
// Equation(s):
// \Mux29~18_combout  = (dcifimemload_22 & ((\Mux29~17_combout  & (\regs[15][2]~q )) # (!\Mux29~17_combout  & ((\regs[14][2]~q ))))) # (!dcifimemload_22 & (\Mux29~17_combout ))

	.dataa(dcifimemload_22),
	.datab(\Mux29~17_combout ),
	.datac(\regs[15][2]~q ),
	.datad(\regs[14][2]~q ),
	.cin(gnd),
	.combout(\Mux29~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~18 .lut_mask = 16'hE6C4;
defparam \Mux29~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N15
dffeas \regs[5][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][2] .is_wysiwyg = "true";
defparam \regs[5][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (dcifimemload_21 & (((\regs[5][2]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][2]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][2]~q ),
	.datac(\regs[5][2]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hAAE4;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N20
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (dcifimemload_22 & ((\Mux29~10_combout  & (\regs[7][2]~q )) # (!\Mux29~10_combout  & ((\regs[6][2]~q ))))) # (!dcifimemload_22 & (((\Mux29~10_combout ))))

	.dataa(\regs[7][2]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[6][2]~q ),
	.datad(\Mux29~10_combout ),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'hBBC0;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N27
dffeas \regs[1][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][2] .is_wysiwyg = "true";
defparam \regs[1][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N26
cycloneive_lcell_comb \Mux29~14 (
// Equation(s):
// \Mux29~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\regs[3][2]~q )) # (!dcifimemload_22 & ((\regs[1][2]~q )))))

	.dataa(dcifimemload_21),
	.datab(\regs[3][2]~q ),
	.datac(\regs[1][2]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux29~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~14 .lut_mask = 16'h88A0;
defparam \Mux29~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N18
cycloneive_lcell_comb \Mux29~15 (
// Equation(s):
// \Mux29~15_combout  = (\Mux29~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][2]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[2][2]~q ),
	.datad(\Mux29~14_combout ),
	.cin(gnd),
	.combout(\Mux29~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~15 .lut_mask = 16'hFF20;
defparam \Mux29~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N23
dffeas \regs[8][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~62_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][2] .is_wysiwyg = "true";
defparam \regs[8][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N22
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// \Mux29~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\regs[10][2]~q )) # (!dcifimemload_22 & ((\regs[8][2]~q )))))

	.dataa(\regs[10][2]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[8][2]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux29~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hEE30;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N16
cycloneive_lcell_comb \Mux29~13 (
// Equation(s):
// \Mux29~13_combout  = (dcifimemload_21 & ((\Mux29~12_combout  & ((\regs[11][2]~q ))) # (!\Mux29~12_combout  & (\regs[9][2]~q )))) # (!dcifimemload_21 & (((\Mux29~12_combout ))))

	.dataa(\regs[9][2]~q ),
	.datab(\regs[11][2]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux29~12_combout ),
	.cin(gnd),
	.combout(\Mux29~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~13 .lut_mask = 16'hCFA0;
defparam \Mux29~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N2
cycloneive_lcell_comb \Mux29~16 (
// Equation(s):
// \Mux29~16_combout  = (dcifimemload_24 & (((dcifimemload_23) # (\Mux29~13_combout )))) # (!dcifimemload_24 & (\Mux29~15_combout  & (!dcifimemload_23)))

	.dataa(dcifimemload_24),
	.datab(\Mux29~15_combout ),
	.datac(dcifimemload_23),
	.datad(\Mux29~13_combout ),
	.cin(gnd),
	.combout(\Mux29~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~16 .lut_mask = 16'hAEA4;
defparam \Mux29~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N0
cycloneive_lcell_comb \Mux29~19 (
// Equation(s):
// \Mux29~19_combout  = (dcifimemload_23 & ((\Mux29~16_combout  & (\Mux29~18_combout )) # (!\Mux29~16_combout  & ((\Mux29~11_combout ))))) # (!dcifimemload_23 & (((\Mux29~16_combout ))))

	.dataa(\Mux29~18_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux29~11_combout ),
	.datad(\Mux29~16_combout ),
	.cin(gnd),
	.combout(\Mux29~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~19 .lut_mask = 16'hBBC0;
defparam \Mux29~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y37_N29
dffeas \regs[16][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][1] .is_wysiwyg = "true";
defparam \regs[16][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N28
cycloneive_lcell_comb \Mux62~4 (
// Equation(s):
// \Mux62~4_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[20][1]~q )) # (!dcifimemload_18 & ((\regs[16][1]~q )))))

	.dataa(dcifimemload_19),
	.datab(\regs[20][1]~q ),
	.datac(\regs[16][1]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux62~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~4 .lut_mask = 16'hEE50;
defparam \Mux62~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N22
cycloneive_lcell_comb \Mux62~5 (
// Equation(s):
// \Mux62~5_combout  = (dcifimemload_19 & ((\Mux62~4_combout  & ((\regs[28][1]~q ))) # (!\Mux62~4_combout  & (\regs[24][1]~q )))) # (!dcifimemload_19 & (((\Mux62~4_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[24][1]~q ),
	.datac(\regs[28][1]~q ),
	.datad(\Mux62~4_combout ),
	.cin(gnd),
	.combout(\Mux62~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~5 .lut_mask = 16'hF588;
defparam \Mux62~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N31
dffeas \regs[30][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][1] .is_wysiwyg = "true";
defparam \regs[30][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N24
cycloneive_lcell_comb \Mux62~2 (
// Equation(s):
// \Mux62~2_combout  = (dcifimemload_18 & ((\regs[22][1]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\regs[18][1]~q  & !dcifimemload_19))))

	.dataa(\regs[22][1]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[18][1]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~2 .lut_mask = 16'hCCB8;
defparam \Mux62~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N30
cycloneive_lcell_comb \Mux62~3 (
// Equation(s):
// \Mux62~3_combout  = (dcifimemload_19 & ((\Mux62~2_combout  & ((\regs[30][1]~q ))) # (!\Mux62~2_combout  & (\regs[26][1]~q )))) # (!dcifimemload_19 & (((\Mux62~2_combout ))))

	.dataa(\regs[26][1]~q ),
	.datab(dcifimemload_19),
	.datac(\regs[30][1]~q ),
	.datad(\Mux62~2_combout ),
	.cin(gnd),
	.combout(\Mux62~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~3 .lut_mask = 16'hF388;
defparam \Mux62~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N20
cycloneive_lcell_comb \Mux62~6 (
// Equation(s):
// \Mux62~6_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux62~3_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux62~5_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux62~5_combout ),
	.datad(\Mux62~3_combout ),
	.cin(gnd),
	.combout(\Mux62~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~6 .lut_mask = 16'hBA98;
defparam \Mux62~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N23
dffeas \regs[17][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][1] .is_wysiwyg = "true";
defparam \regs[17][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N22
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (dcifimemload_19 & ((\regs[25][1]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\regs[17][1]~q  & !dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\regs[25][1]~q ),
	.datac(\regs[17][1]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hAAD8;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N30
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (dcifimemload_18 & ((\Mux62~0_combout  & ((\regs[29][1]~q ))) # (!\Mux62~0_combout  & (\regs[21][1]~q )))) # (!dcifimemload_18 & (((\Mux62~0_combout ))))

	.dataa(\regs[21][1]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[29][1]~q ),
	.datad(\Mux62~0_combout ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hF388;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N12
cycloneive_lcell_comb \regs[23][1]~feeder (
// Equation(s):
// \regs[23][1]~feeder_combout  = \regs~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~7_combout ),
	.cin(gnd),
	.combout(\regs[23][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][1]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N13
dffeas \regs[23][1] (
	.clk(CLK),
	.d(\regs[23][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][1] .is_wysiwyg = "true";
defparam \regs[23][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N12
cycloneive_lcell_comb \Mux62~7 (
// Equation(s):
// \Mux62~7_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[27][1]~q )) # (!dcifimemload_19 & ((\regs[19][1]~q )))))

	.dataa(\regs[27][1]~q ),
	.datab(\regs[19][1]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux62~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~7 .lut_mask = 16'hFA0C;
defparam \Mux62~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N2
cycloneive_lcell_comb \Mux62~8 (
// Equation(s):
// \Mux62~8_combout  = (dcifimemload_18 & ((\Mux62~7_combout  & (\regs[31][1]~q )) # (!\Mux62~7_combout  & ((\regs[23][1]~q ))))) # (!dcifimemload_18 & (((\Mux62~7_combout ))))

	.dataa(\regs[31][1]~q ),
	.datab(\regs[23][1]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux62~7_combout ),
	.cin(gnd),
	.combout(\Mux62~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~8 .lut_mask = 16'hAFC0;
defparam \Mux62~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N31
dffeas \regs[4][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][1] .is_wysiwyg = "true";
defparam \regs[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \Mux62~10 (
// Equation(s):
// \Mux62~10_combout  = (dcifimemload_16 & ((\regs[5][1]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\regs[4][1]~q  & !dcifimemload_17))))

	.dataa(\regs[5][1]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[4][1]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux62~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~10 .lut_mask = 16'hCCB8;
defparam \Mux62~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N14
cycloneive_lcell_comb \Mux62~11 (
// Equation(s):
// \Mux62~11_combout  = (dcifimemload_17 & ((\Mux62~10_combout  & (\regs[7][1]~q )) # (!\Mux62~10_combout  & ((\regs[6][1]~q ))))) # (!dcifimemload_17 & (\Mux62~10_combout ))

	.dataa(dcifimemload_17),
	.datab(\Mux62~10_combout ),
	.datac(\regs[7][1]~q ),
	.datad(\regs[6][1]~q ),
	.cin(gnd),
	.combout(\Mux62~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~11 .lut_mask = 16'hE6C4;
defparam \Mux62~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N24
cycloneive_lcell_comb \Mux62~17 (
// Equation(s):
// \Mux62~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][1]~q )) # (!dcifimemload_16 & ((\regs[12][1]~q )))))

	.dataa(dcifimemload_17),
	.datab(\regs[13][1]~q ),
	.datac(\regs[12][1]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux62~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~17 .lut_mask = 16'hEE50;
defparam \Mux62~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N18
cycloneive_lcell_comb \Mux62~18 (
// Equation(s):
// \Mux62~18_combout  = (\Mux62~17_combout  & (((\regs[15][1]~q ) # (!dcifimemload_17)))) # (!\Mux62~17_combout  & (\regs[14][1]~q  & ((dcifimemload_17))))

	.dataa(\regs[14][1]~q ),
	.datab(\Mux62~17_combout ),
	.datac(\regs[15][1]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux62~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~18 .lut_mask = 16'hE2CC;
defparam \Mux62~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N15
dffeas \regs[11][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][1] .is_wysiwyg = "true";
defparam \regs[11][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N29
dffeas \regs[8][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][1] .is_wysiwyg = "true";
defparam \regs[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N28
cycloneive_lcell_comb \Mux62~12 (
// Equation(s):
// \Mux62~12_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][1]~q )) # (!dcifimemload_17 & ((\regs[8][1]~q )))))

	.dataa(\regs[10][1]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[8][1]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux62~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~12 .lut_mask = 16'hEE30;
defparam \Mux62~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N14
cycloneive_lcell_comb \Mux62~13 (
// Equation(s):
// \Mux62~13_combout  = (dcifimemload_16 & ((\Mux62~12_combout  & ((\regs[11][1]~q ))) # (!\Mux62~12_combout  & (\regs[9][1]~q )))) # (!dcifimemload_16 & (((\Mux62~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][1]~q ),
	.datac(\regs[11][1]~q ),
	.datad(\Mux62~12_combout ),
	.cin(gnd),
	.combout(\Mux62~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~13 .lut_mask = 16'hF588;
defparam \Mux62~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N13
dffeas \regs[2][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][1] .is_wysiwyg = "true";
defparam \regs[2][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N16
cycloneive_lcell_comb \Mux62~14 (
// Equation(s):
// \Mux62~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\regs[3][1]~q ))) # (!dcifimemload_17 & (\regs[1][1]~q ))))

	.dataa(\regs[1][1]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[3][1]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux62~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~14 .lut_mask = 16'hC088;
defparam \Mux62~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N12
cycloneive_lcell_comb \Mux62~15 (
// Equation(s):
// \Mux62~15_combout  = (\Mux62~14_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \regs[2][1]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\regs[2][1]~q ),
	.datad(\Mux62~14_combout ),
	.cin(gnd),
	.combout(\Mux62~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~15 .lut_mask = 16'hFF40;
defparam \Mux62~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N6
cycloneive_lcell_comb \Mux62~16 (
// Equation(s):
// \Mux62~16_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux62~13_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & ((\Mux62~15_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux62~13_combout ),
	.datad(\Mux62~15_combout ),
	.cin(gnd),
	.combout(\Mux62~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~16 .lut_mask = 16'hB9A8;
defparam \Mux62~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N16
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (dcifimemload_24 & (((\regs[25][0]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[17][0]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[17][0]~q ),
	.datac(\regs[25][0]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hAAE4;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N10
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (\Mux31~0_combout  & (((\regs[29][0]~q ) # (!dcifimemload_23)))) # (!\Mux31~0_combout  & (\regs[21][0]~q  & ((dcifimemload_23))))

	.dataa(\regs[21][0]~q ),
	.datab(\regs[29][0]~q ),
	.datac(\Mux31~0_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hCAF0;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N2
cycloneive_lcell_comb \regs[26][0]~feeder (
// Equation(s):
// \regs[26][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[26][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][0]~feeder .lut_mask = 16'hF0F0;
defparam \regs[26][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N3
dffeas \regs[26][0] (
	.clk(CLK),
	.d(\regs[26][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][0] .is_wysiwyg = "true";
defparam \regs[26][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N2
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[22][0]~q )) # (!dcifimemload_23 & ((\regs[18][0]~q )))))

	.dataa(\regs[22][0]~q ),
	.datab(\regs[18][0]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hFA0C;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N16
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (dcifimemload_24 & ((\Mux31~2_combout  & ((\regs[30][0]~q ))) # (!\Mux31~2_combout  & (\regs[26][0]~q )))) # (!dcifimemload_24 & (((\Mux31~2_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[26][0]~q ),
	.datac(\regs[30][0]~q ),
	.datad(\Mux31~2_combout ),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hF588;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N18
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (dcifimemload_23 & (((\regs[20][0]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\regs[16][0]~q  & ((!dcifimemload_24))))

	.dataa(\regs[16][0]~q ),
	.datab(\regs[20][0]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hF0CA;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N10
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (dcifimemload_24 & ((\Mux31~4_combout  & (\regs[28][0]~q )) # (!\Mux31~4_combout  & ((\regs[24][0]~q ))))) # (!dcifimemload_24 & (((\Mux31~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\regs[28][0]~q ),
	.datac(\regs[24][0]~q ),
	.datad(\Mux31~4_combout ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hDDA0;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N4
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux31~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux31~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux31~3_combout ),
	.datad(\Mux31~5_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hB9A8;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N8
cycloneive_lcell_comb \regs[19][0]~feeder (
// Equation(s):
// \regs[19][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~5_combout ),
	.cin(gnd),
	.combout(\regs[19][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][0]~feeder .lut_mask = 16'hFF00;
defparam \regs[19][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N9
dffeas \regs[19][0] (
	.clk(CLK),
	.d(\regs[19][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][0] .is_wysiwyg = "true";
defparam \regs[19][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N8
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (dcifimemload_24 & (((\regs[27][0]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\regs[19][0]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\regs[19][0]~q ),
	.datac(\regs[27][0]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hAAE4;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N16
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (dcifimemload_23 & ((\Mux31~7_combout  & ((\regs[31][0]~q ))) # (!\Mux31~7_combout  & (\regs[23][0]~q )))) # (!dcifimemload_23 & (((\Mux31~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[23][0]~q ),
	.datac(\regs[31][0]~q ),
	.datad(\Mux31~7_combout ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hF588;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N26
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// \Mux31~9_combout  = (dcifimemload_21 & ((\Mux31~6_combout  & ((\Mux31~8_combout ))) # (!\Mux31~6_combout  & (\Mux31~1_combout )))) # (!dcifimemload_21 & (((\Mux31~6_combout ))))

	.dataa(\Mux31~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux31~6_combout ),
	.datad(\Mux31~8_combout ),
	.cin(gnd),
	.combout(\Mux31~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hF838;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N9
dffeas \regs[6][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][0] .is_wysiwyg = "true";
defparam \regs[6][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N18
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (dcifimemload_21 & (((\regs[5][0]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][0]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\regs[4][0]~q ),
	.datac(\regs[5][0]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hAAE4;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N8
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (dcifimemload_22 & ((\Mux31~10_combout  & (\regs[7][0]~q )) # (!\Mux31~10_combout  & ((\regs[6][0]~q ))))) # (!dcifimemload_22 & (((\Mux31~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[7][0]~q ),
	.datac(\regs[6][0]~q ),
	.datad(\Mux31~10_combout ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'hDDA0;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// \Mux31~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\regs[10][0]~q ))) # (!dcifimemload_22 & (\regs[8][0]~q ))))

	.dataa(dcifimemload_21),
	.datab(\regs[8][0]~q ),
	.datac(\regs[10][0]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux31~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hFA44;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N0
cycloneive_lcell_comb \Mux31~13 (
// Equation(s):
// \Mux31~13_combout  = (dcifimemload_21 & ((\Mux31~12_combout  & (\regs[11][0]~q )) # (!\Mux31~12_combout  & ((\regs[9][0]~q ))))) # (!dcifimemload_21 & (((\Mux31~12_combout ))))

	.dataa(\regs[11][0]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[9][0]~q ),
	.datad(\Mux31~12_combout ),
	.cin(gnd),
	.combout(\Mux31~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~13 .lut_mask = 16'hBBC0;
defparam \Mux31~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N11
dffeas \regs[2][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][0] .is_wysiwyg = "true";
defparam \regs[2][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N28
cycloneive_lcell_comb \Mux31~14 (
// Equation(s):
// \Mux31~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][0]~q ))) # (!dcifimemload_22 & (\regs[1][0]~q ))))

	.dataa(dcifimemload_22),
	.datab(\regs[1][0]~q ),
	.datac(dcifimemload_21),
	.datad(\regs[3][0]~q ),
	.cin(gnd),
	.combout(\Mux31~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~14 .lut_mask = 16'hE040;
defparam \Mux31~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N10
cycloneive_lcell_comb \Mux31~15 (
// Equation(s):
// \Mux31~15_combout  = (\Mux31~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \regs[2][0]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[2][0]~q ),
	.datad(\Mux31~14_combout ),
	.cin(gnd),
	.combout(\Mux31~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~15 .lut_mask = 16'hFF20;
defparam \Mux31~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N22
cycloneive_lcell_comb \Mux31~16 (
// Equation(s):
// \Mux31~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & (\Mux31~13_combout )) # (!dcifimemload_24 & ((\Mux31~15_combout )))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux31~13_combout ),
	.datad(\Mux31~15_combout ),
	.cin(gnd),
	.combout(\Mux31~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~16 .lut_mask = 16'hD9C8;
defparam \Mux31~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N12
cycloneive_lcell_comb \regs[13][0]~feeder (
// Equation(s):
// \regs[13][0]~feeder_combout  = \regs~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~5_combout ),
	.cin(gnd),
	.combout(\regs[13][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][0]~feeder .lut_mask = 16'hFF00;
defparam \regs[13][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N13
dffeas \regs[13][0] (
	.clk(CLK),
	.d(\regs[13][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][0] .is_wysiwyg = "true";
defparam \regs[13][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N14
cycloneive_lcell_comb \Mux31~17 (
// Equation(s):
// \Mux31~17_combout  = (dcifimemload_21 & (((\regs[13][0]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[12][0]~q  & ((!dcifimemload_22))))

	.dataa(\regs[12][0]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[13][0]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux31~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~17 .lut_mask = 16'hCCE2;
defparam \Mux31~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N26
cycloneive_lcell_comb \Mux31~18 (
// Equation(s):
// \Mux31~18_combout  = (dcifimemload_22 & ((\Mux31~17_combout  & (\regs[15][0]~q )) # (!\Mux31~17_combout  & ((\regs[14][0]~q ))))) # (!dcifimemload_22 & (((\Mux31~17_combout ))))

	.dataa(\regs[15][0]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[14][0]~q ),
	.datad(\Mux31~17_combout ),
	.cin(gnd),
	.combout(\Mux31~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~18 .lut_mask = 16'hBBC0;
defparam \Mux31~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N20
cycloneive_lcell_comb \Mux31~19 (
// Equation(s):
// \Mux31~19_combout  = (dcifimemload_23 & ((\Mux31~16_combout  & ((\Mux31~18_combout ))) # (!\Mux31~16_combout  & (\Mux31~11_combout )))) # (!dcifimemload_23 & (((\Mux31~16_combout ))))

	.dataa(\Mux31~11_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux31~16_combout ),
	.datad(\Mux31~18_combout ),
	.cin(gnd),
	.combout(\Mux31~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~19 .lut_mask = 16'hF838;
defparam \Mux31~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N20
cycloneive_lcell_comb \regs~63 (
// Equation(s):
// \regs~63_combout  = (\Selector0~1_combout  & !\Equal0~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector01),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\regs~63_combout ),
	.cout());
// synopsys translate_off
defparam \regs~63 .lut_mask = 16'h00F0;
defparam \regs~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N5
dffeas \regs[14][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][31] .is_wysiwyg = "true";
defparam \regs[14][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N19
dffeas \regs[15][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][31] .is_wysiwyg = "true";
defparam \regs[15][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y44_N27
dffeas \regs[12][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][31] .is_wysiwyg = "true";
defparam \regs[12][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N26
cycloneive_lcell_comb \Mux32~7 (
// Equation(s):
// \Mux32~7_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\regs[13][31]~q )) # (!dcifimemload_16 & ((\regs[12][31]~q )))))

	.dataa(\regs[13][31]~q ),
	.datab(dcifimemload_17),
	.datac(\regs[12][31]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux32~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~7 .lut_mask = 16'hEE30;
defparam \Mux32~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N18
cycloneive_lcell_comb \Mux32~8 (
// Equation(s):
// \Mux32~8_combout  = (dcifimemload_17 & ((\Mux32~7_combout  & ((\regs[15][31]~q ))) # (!\Mux32~7_combout  & (\regs[14][31]~q )))) # (!dcifimemload_17 & (((\Mux32~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\regs[14][31]~q ),
	.datac(\regs[15][31]~q ),
	.datad(\Mux32~7_combout ),
	.cin(gnd),
	.combout(\Mux32~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~8 .lut_mask = 16'hF588;
defparam \Mux32~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N31
dffeas \regs[7][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][31] .is_wysiwyg = "true";
defparam \regs[7][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N28
cycloneive_lcell_comb \regs[6][31]~feeder (
// Equation(s):
// \regs[6][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~63_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[6][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][31]~feeder .lut_mask = 16'hF0F0;
defparam \regs[6][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N29
dffeas \regs[6][31] (
	.clk(CLK),
	.d(\regs[6][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][31] .is_wysiwyg = "true";
defparam \regs[6][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N20
cycloneive_lcell_comb \regs[5][31]~feeder (
// Equation(s):
// \regs[5][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~63_combout ),
	.cin(gnd),
	.combout(\regs[5][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[5][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N21
dffeas \regs[5][31] (
	.clk(CLK),
	.d(\regs[5][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][31] .is_wysiwyg = "true";
defparam \regs[5][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N0
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\regs[5][31]~q ))) # (!dcifimemload_16 & (\regs[4][31]~q ))))

	.dataa(\regs[4][31]~q ),
	.datab(\regs[5][31]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hFC0A;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N12
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (dcifimemload_17 & ((\Mux32~0_combout  & (\regs[7][31]~q )) # (!\Mux32~0_combout  & ((\regs[6][31]~q ))))) # (!dcifimemload_17 & (((\Mux32~0_combout ))))

	.dataa(\regs[7][31]~q ),
	.datab(\regs[6][31]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux32~0_combout ),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hAFC0;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N11
dffeas \regs[2][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][31] .is_wysiwyg = "true";
defparam \regs[2][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y42_N29
dffeas \regs[1][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][31] .is_wysiwyg = "true";
defparam \regs[1][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N28
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\regs[3][31]~q )) # (!dcifimemload_17 & ((\regs[1][31]~q )))))

	.dataa(\regs[3][31]~q ),
	.datab(dcifimemload_16),
	.datac(\regs[1][31]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'h88C0;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N10
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (\Mux32~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \regs[2][31]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\regs[2][31]~q ),
	.datad(\Mux32~4_combout ),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'hFF20;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N1
dffeas \regs[9][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][31] .is_wysiwyg = "true";
defparam \regs[9][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N23
dffeas \regs[11][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][31] .is_wysiwyg = "true";
defparam \regs[11][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N3
dffeas \regs[10][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][31] .is_wysiwyg = "true";
defparam \regs[10][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N1
dffeas \regs[8][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][31] .is_wysiwyg = "true";
defparam \regs[8][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N0
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\regs[10][31]~q )) # (!dcifimemload_17 & ((\regs[8][31]~q )))))

	.dataa(dcifimemload_16),
	.datab(\regs[10][31]~q ),
	.datac(\regs[8][31]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'hEE50;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N22
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (dcifimemload_16 & ((\Mux32~2_combout  & ((\regs[11][31]~q ))) # (!\Mux32~2_combout  & (\regs[9][31]~q )))) # (!dcifimemload_16 & (((\Mux32~2_combout ))))

	.dataa(dcifimemload_16),
	.datab(\regs[9][31]~q ),
	.datac(\regs[11][31]~q ),
	.datad(\Mux32~2_combout ),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hF588;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N2
cycloneive_lcell_comb \Mux32~6 (
// Equation(s):
// \Mux32~6_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux32~3_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & (\Mux32~5_combout )))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux32~5_combout ),
	.datad(\Mux32~3_combout ),
	.cin(gnd),
	.combout(\Mux32~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~6 .lut_mask = 16'hBA98;
defparam \Mux32~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N26
cycloneive_lcell_comb \regs[31][31]~feeder (
// Equation(s):
// \regs[31][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~63_combout ),
	.cin(gnd),
	.combout(\regs[31][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[31][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N27
dffeas \regs[31][31] (
	.clk(CLK),
	.d(\regs[31][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][31] .is_wysiwyg = "true";
defparam \regs[31][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N5
dffeas \regs[23][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][31] .is_wysiwyg = "true";
defparam \regs[23][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y44_N20
cycloneive_lcell_comb \regs[19][31]~feeder (
// Equation(s):
// \regs[19][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~63_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[19][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][31]~feeder .lut_mask = 16'hF0F0;
defparam \regs[19][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y44_N21
dffeas \regs[19][31] (
	.clk(CLK),
	.d(\regs[19][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][31] .is_wysiwyg = "true";
defparam \regs[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N20
cycloneive_lcell_comb \Mux32~17 (
// Equation(s):
// \Mux32~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[27][31]~q )) # (!dcifimemload_19 & ((\regs[19][31]~q )))))

	.dataa(\regs[27][31]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[19][31]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux32~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~17 .lut_mask = 16'hEE30;
defparam \Mux32~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N2
cycloneive_lcell_comb \Mux32~18 (
// Equation(s):
// \Mux32~18_combout  = (dcifimemload_18 & ((\Mux32~17_combout  & (\regs[31][31]~q )) # (!\Mux32~17_combout  & ((\regs[23][31]~q ))))) # (!dcifimemload_18 & (((\Mux32~17_combout ))))

	.dataa(\regs[31][31]~q ),
	.datab(dcifimemload_18),
	.datac(\regs[23][31]~q ),
	.datad(\Mux32~17_combout ),
	.cin(gnd),
	.combout(\Mux32~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~18 .lut_mask = 16'hBBC0;
defparam \Mux32~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N18
cycloneive_lcell_comb \regs[29][31]~feeder (
// Equation(s):
// \regs[29][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~63_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[29][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][31]~feeder .lut_mask = 16'hF0F0;
defparam \regs[29][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N19
dffeas \regs[29][31] (
	.clk(CLK),
	.d(\regs[29][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][31] .is_wysiwyg = "true";
defparam \regs[29][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N16
cycloneive_lcell_comb \regs[21][31]~feeder (
// Equation(s):
// \regs[21][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\regs~63_combout ),
	.cin(gnd),
	.combout(\regs[21][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[21][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N17
dffeas \regs[21][31] (
	.clk(CLK),
	.d(\regs[21][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][31] .is_wysiwyg = "true";
defparam \regs[21][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N16
cycloneive_lcell_comb \regs[17][31]~feeder (
// Equation(s):
// \regs[17][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~63_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[17][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][31]~feeder .lut_mask = 16'hF0F0;
defparam \regs[17][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N17
dffeas \regs[17][31] (
	.clk(CLK),
	.d(\regs[17][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][31] .is_wysiwyg = "true";
defparam \regs[17][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N12
cycloneive_lcell_comb \Mux32~10 (
// Equation(s):
// \Mux32~10_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\regs[25][31]~q )) # (!dcifimemload_19 & ((\regs[17][31]~q )))))

	.dataa(\regs[25][31]~q ),
	.datab(\regs[17][31]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux32~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~10 .lut_mask = 16'hFA0C;
defparam \Mux32~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N18
cycloneive_lcell_comb \Mux32~11 (
// Equation(s):
// \Mux32~11_combout  = (dcifimemload_18 & ((\Mux32~10_combout  & (\regs[29][31]~q )) # (!\Mux32~10_combout  & ((\regs[21][31]~q ))))) # (!dcifimemload_18 & (((\Mux32~10_combout ))))

	.dataa(\regs[29][31]~q ),
	.datab(\regs[21][31]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux32~10_combout ),
	.cin(gnd),
	.combout(\Mux32~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~11 .lut_mask = 16'hAFC0;
defparam \Mux32~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N19
dffeas \regs[28][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][31] .is_wysiwyg = "true";
defparam \regs[28][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N5
dffeas \regs[24][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][31] .is_wysiwyg = "true";
defparam \regs[24][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N7
dffeas \regs[20][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][31] .is_wysiwyg = "true";
defparam \regs[20][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N29
dffeas \regs[16][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][31] .is_wysiwyg = "true";
defparam \regs[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N6
cycloneive_lcell_comb \Mux32~14 (
// Equation(s):
// \Mux32~14_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & (\regs[20][31]~q )) # (!dcifimemload_18 & ((\regs[16][31]~q )))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\regs[20][31]~q ),
	.datad(\regs[16][31]~q ),
	.cin(gnd),
	.combout(\Mux32~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~14 .lut_mask = 16'hD9C8;
defparam \Mux32~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N4
cycloneive_lcell_comb \Mux32~15 (
// Equation(s):
// \Mux32~15_combout  = (dcifimemload_19 & ((\Mux32~14_combout  & (\regs[28][31]~q )) # (!\Mux32~14_combout  & ((\regs[24][31]~q ))))) # (!dcifimemload_19 & (((\Mux32~14_combout ))))

	.dataa(dcifimemload_19),
	.datab(\regs[28][31]~q ),
	.datac(\regs[24][31]~q ),
	.datad(\Mux32~14_combout ),
	.cin(gnd),
	.combout(\Mux32~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~15 .lut_mask = 16'hDDA0;
defparam \Mux32~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N8
cycloneive_lcell_comb \regs[26][31]~feeder (
// Equation(s):
// \regs[26][31]~feeder_combout  = \regs~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\regs~63_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[26][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[26][31]~feeder .lut_mask = 16'hF0F0;
defparam \regs[26][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N9
dffeas \regs[26][31] (
	.clk(CLK),
	.d(\regs[26][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][31] .is_wysiwyg = "true";
defparam \regs[26][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N9
dffeas \regs[18][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][31] .is_wysiwyg = "true";
defparam \regs[18][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N19
dffeas \regs[22][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][31] .is_wysiwyg = "true";
defparam \regs[22][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N18
cycloneive_lcell_comb \Mux32~12 (
// Equation(s):
// \Mux32~12_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\regs[22][31]~q ))) # (!dcifimemload_18 & (\regs[18][31]~q ))))

	.dataa(dcifimemload_19),
	.datab(\regs[18][31]~q ),
	.datac(\regs[22][31]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux32~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~12 .lut_mask = 16'hFA44;
defparam \Mux32~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N16
cycloneive_lcell_comb \Mux32~13 (
// Equation(s):
// \Mux32~13_combout  = (dcifimemload_19 & ((\Mux32~12_combout  & (\regs[30][31]~q )) # (!\Mux32~12_combout  & ((\regs[26][31]~q ))))) # (!dcifimemload_19 & (((\Mux32~12_combout ))))

	.dataa(\regs[30][31]~q ),
	.datab(\regs[26][31]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux32~12_combout ),
	.cin(gnd),
	.combout(\Mux32~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~13 .lut_mask = 16'hAFC0;
defparam \Mux32~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N12
cycloneive_lcell_comb \Mux32~16 (
// Equation(s):
// \Mux32~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux32~13_combout ))) # (!dcifimemload_17 & (\Mux32~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux32~15_combout ),
	.datad(\Mux32~13_combout ),
	.cin(gnd),
	.combout(\Mux32~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~16 .lut_mask = 16'hDC98;
defparam \Mux32~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y44_N25
dffeas \regs[13][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][31] .is_wysiwyg = "true";
defparam \regs[13][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y44_N24
cycloneive_lcell_comb \Mux0~17 (
// Equation(s):
// \Mux0~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\regs[13][31]~q ))) # (!dcifimemload_21 & (\regs[12][31]~q ))))

	.dataa(\regs[12][31]~q ),
	.datab(dcifimemload_22),
	.datac(\regs[13][31]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~17 .lut_mask = 16'hFC22;
defparam \Mux0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N4
cycloneive_lcell_comb \Mux0~18 (
// Equation(s):
// \Mux0~18_combout  = (dcifimemload_22 & ((\Mux0~17_combout  & (\regs[15][31]~q )) # (!\Mux0~17_combout  & ((\regs[14][31]~q ))))) # (!dcifimemload_22 & (((\Mux0~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[15][31]~q ),
	.datac(\regs[14][31]~q ),
	.datad(\Mux0~17_combout ),
	.cin(gnd),
	.combout(\Mux0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~18 .lut_mask = 16'hDDA0;
defparam \Mux0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N2
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\regs[10][31]~q )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\regs[8][31]~q ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\regs[10][31]~q ),
	.datad(\regs[8][31]~q ),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'hB9A8;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N0
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (dcifimemload_21 & ((\Mux0~10_combout  & (\regs[11][31]~q )) # (!\Mux0~10_combout  & ((\regs[9][31]~q ))))) # (!dcifimemload_21 & (((\Mux0~10_combout ))))

	.dataa(\regs[11][31]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[9][31]~q ),
	.datad(\Mux0~10_combout ),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hBBC0;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N9
dffeas \regs[3][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][31] .is_wysiwyg = "true";
defparam \regs[3][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N8
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// \Mux0~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\regs[3][31]~q ))) # (!dcifimemload_22 & (\regs[1][31]~q ))))

	.dataa(\regs[1][31]~q ),
	.datab(dcifimemload_21),
	.datac(\regs[3][31]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'hC088;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N30
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// \Mux0~15_combout  = (\Mux0~14_combout ) # ((\regs[2][31]~q  & (!dcifimemload_21 & dcifimemload_22)))

	.dataa(\regs[2][31]~q ),
	.datab(dcifimemload_21),
	.datac(\Mux0~14_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hF2F0;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N18
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (dcifimemload_21 & (((\regs[5][31]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\regs[4][31]~q  & ((!dcifimemload_22))))

	.dataa(\regs[4][31]~q ),
	.datab(\regs[5][31]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hF0CA;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N30
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// \Mux0~13_combout  = (dcifimemload_22 & ((\Mux0~12_combout  & ((\regs[7][31]~q ))) # (!\Mux0~12_combout  & (\regs[6][31]~q )))) # (!dcifimemload_22 & (((\Mux0~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\regs[6][31]~q ),
	.datac(\regs[7][31]~q ),
	.datad(\Mux0~12_combout ),
	.cin(gnd),
	.combout(\Mux0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hF588;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N24
cycloneive_lcell_comb \Mux0~16 (
// Equation(s):
// \Mux0~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux0~13_combout ))) # (!dcifimemload_23 & (\Mux0~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux0~15_combout ),
	.datad(\Mux0~13_combout ),
	.cin(gnd),
	.combout(\Mux0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~16 .lut_mask = 16'hDC98;
defparam \Mux0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N22
cycloneive_lcell_comb \Mux0~19 (
// Equation(s):
// \Mux0~19_combout  = (dcifimemload_24 & ((\Mux0~16_combout  & (\Mux0~18_combout )) # (!\Mux0~16_combout  & ((\Mux0~11_combout ))))) # (!dcifimemload_24 & (((\Mux0~16_combout ))))

	.dataa(\Mux0~18_combout ),
	.datab(\Mux0~11_combout ),
	.datac(dcifimemload_24),
	.datad(\Mux0~16_combout ),
	.cin(gnd),
	.combout(\Mux0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~19 .lut_mask = 16'hAFC0;
defparam \Mux0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N28
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\regs[21][31]~q )) # (!dcifimemload_23 & ((\regs[17][31]~q )))))

	.dataa(\regs[21][31]~q ),
	.datab(\regs[17][31]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hFA0C;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N2
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (dcifimemload_24 & ((\Mux0~0_combout  & ((\regs[29][31]~q ))) # (!\Mux0~0_combout  & (\regs[25][31]~q )))) # (!dcifimemload_24 & (((\Mux0~0_combout ))))

	.dataa(\regs[25][31]~q ),
	.datab(\regs[29][31]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hCFA0;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N4
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (dcifimemload_23 & ((\regs[23][31]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\regs[19][31]~q  & !dcifimemload_24))))

	.dataa(\regs[23][31]~q ),
	.datab(\regs[19][31]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hF0AC;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N2
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (\Mux0~7_combout  & (((\regs[31][31]~q ) # (!dcifimemload_24)))) # (!\Mux0~7_combout  & (\regs[27][31]~q  & ((dcifimemload_24))))

	.dataa(\regs[27][31]~q ),
	.datab(\Mux0~7_combout ),
	.datac(\regs[31][31]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'hE2CC;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N28
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & ((\regs[24][31]~q ))) # (!dcifimemload_24 & (\regs[16][31]~q ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\regs[16][31]~q ),
	.datad(\regs[24][31]~q ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'hDC98;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N18
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (dcifimemload_23 & ((\Mux0~4_combout  & ((\regs[28][31]~q ))) # (!\Mux0~4_combout  & (\regs[20][31]~q )))) # (!dcifimemload_23 & (((\Mux0~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\regs[20][31]~q ),
	.datac(\regs[28][31]~q ),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hF588;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N3
dffeas \regs[30][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\regs~63_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][31] .is_wysiwyg = "true";
defparam \regs[30][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N8
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\regs[26][31]~q )) # (!dcifimemload_24 & ((\regs[18][31]~q )))))

	.dataa(\regs[26][31]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[18][31]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hEE30;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N2
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (dcifimemload_23 & ((\Mux0~2_combout  & ((\regs[30][31]~q ))) # (!\Mux0~2_combout  & (\regs[22][31]~q )))) # (!dcifimemload_23 & (((\Mux0~2_combout ))))

	.dataa(\regs[22][31]~q ),
	.datab(dcifimemload_23),
	.datac(\regs[30][31]~q ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'hF388;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N28
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux0~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux0~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux0~5_combout ),
	.datad(\Mux0~3_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hBA98;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N14
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// \Mux0~9_combout  = (dcifimemload_21 & ((\Mux0~6_combout  & ((\Mux0~8_combout ))) # (!\Mux0~6_combout  & (\Mux0~1_combout )))) # (!dcifimemload_21 & (((\Mux0~6_combout ))))

	.dataa(\Mux0~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux0~8_combout ),
	.datad(\Mux0~6_combout ),
	.cin(gnd),
	.combout(\Mux0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hF388;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module request_unit (
	dpifhalt,
	ruifdWEN_r,
	ruifdREN_r,
	always1,
	dcifimemload_26,
	dcifimemload_27,
	dcifimemload_28,
	dcifimemload_29,
	dcifimemload_30,
	dcifimemload_31,
	nxtwen,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	dpifhalt;
output 	ruifdWEN_r;
output 	ruifdREN_r;
input 	always1;
input 	dcifimemload_26;
input 	dcifimemload_27;
input 	dcifimemload_28;
input 	dcifimemload_29;
input 	dcifimemload_30;
input 	dcifimemload_31;
output 	nxtwen;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \nxtwen~6_combout ;
wire \nxtwen~5_combout ;
wire \nxtwen~7_combout ;
wire \nxtren~0_combout ;


// Location: FF_X54_Y37_N9
dffeas \ruif.dWEN_r (
	.clk(CPUCLK),
	.d(\nxtwen~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nxtwen~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ruifdWEN_r),
	.prn(vcc));
// synopsys translate_off
defparam \ruif.dWEN_r .is_wysiwyg = "true";
defparam \ruif.dWEN_r .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N27
dffeas \ruif.dREN_r (
	.clk(CPUCLK),
	.d(\nxtren~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nxtwen~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ruifdREN_r),
	.prn(vcc));
// synopsys translate_off
defparam \ruif.dREN_r .is_wysiwyg = "true";
defparam \ruif.dREN_r .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N16
cycloneive_lcell_comb \nxtwen~4 (
// Equation(s):
// nxtwen = (dcifimemload_26 & (dcifimemload_27 & (dcifimemload_31 & !dcifimemload_28)))

	.dataa(dcifimemload_26),
	.datab(dcifimemload_27),
	.datac(dcifimemload_31),
	.datad(dcifimemload_28),
	.cin(gnd),
	.combout(nxtwen),
	.cout());
// synopsys translate_off
defparam \nxtwen~4 .lut_mask = 16'h0080;
defparam \nxtwen~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N28
cycloneive_lcell_comb \nxtwen~6 (
// Equation(s):
// \nxtwen~6_combout  = (!dpifhalt & (((!ruifdWEN_r & !ruifdREN_r)) # (!always1)))

	.dataa(ruifdWEN_r),
	.datab(ruifdREN_r),
	.datac(dpifhalt),
	.datad(always1),
	.cin(gnd),
	.combout(\nxtwen~6_combout ),
	.cout());
// synopsys translate_off
defparam \nxtwen~6 .lut_mask = 16'h010F;
defparam \nxtwen~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N8
cycloneive_lcell_comb \nxtwen~5 (
// Equation(s):
// \nxtwen~5_combout  = (!dcifimemload_30 & (\nxtwen~6_combout  & (dcifimemload_29 & nxtwen)))

	.dataa(dcifimemload_30),
	.datab(\nxtwen~6_combout ),
	.datac(dcifimemload_29),
	.datad(nxtwen),
	.cin(gnd),
	.combout(\nxtwen~5_combout ),
	.cout());
// synopsys translate_off
defparam \nxtwen~5 .lut_mask = 16'h4000;
defparam \nxtwen~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N30
cycloneive_lcell_comb \nxtwen~7 (
// Equation(s):
// \nxtwen~7_combout  = (always1 & ((ruifdREN_r) # ((ruifdWEN_r) # (!dpifhalt))))

	.dataa(ruifdREN_r),
	.datab(always1),
	.datac(ruifdWEN_r),
	.datad(dpifhalt),
	.cin(gnd),
	.combout(\nxtwen~7_combout ),
	.cout());
// synopsys translate_off
defparam \nxtwen~7 .lut_mask = 16'hC8CC;
defparam \nxtwen~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N26
cycloneive_lcell_comb \nxtren~0 (
// Equation(s):
// \nxtren~0_combout  = (!dcifimemload_30 & (\nxtwen~6_combout  & (!dcifimemload_29 & nxtwen)))

	.dataa(dcifimemload_30),
	.datab(\nxtwen~6_combout ),
	.datac(dcifimemload_29),
	.datad(nxtwen),
	.cin(gnd),
	.combout(\nxtren~0_combout ),
	.cout());
// synopsys translate_off
defparam \nxtren~0 .lut_mask = 16'h0400;
defparam \nxtren~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module memory_control (
	LessThan1,
	ruifdWEN_r,
	ruifdREN_r,
	always0,
	always01,
	always02,
	ccifiwait_0,
	ccifiwait_01,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	LessThan1;
input 	ruifdWEN_r;
input 	ruifdREN_r;
input 	always0;
input 	always01;
input 	always02;
output 	ccifiwait_0;
output 	ccifiwait_01;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \ccif.iwait[0]~1_combout ;


// Location: LCCOMB_X54_Y37_N24
cycloneive_lcell_comb \ccif.iwait[0]~0 (
// Equation(s):
// ccifiwait_0 = (!ruifdWEN_r & !ruifdREN_r)

	.dataa(gnd),
	.datab(ruifdWEN_r),
	.datac(ruifdREN_r),
	.datad(gnd),
	.cin(gnd),
	.combout(ccifiwait_0),
	.cout());
// synopsys translate_off
defparam \ccif.iwait[0]~0 .lut_mask = 16'h0303;
defparam \ccif.iwait[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N2
cycloneive_lcell_comb \ccif.iwait[0] (
// Equation(s):
// ccifiwait_01 = (\ccif.iwait[0]~1_combout ) # ((\nRST~input_o  & ((!always02) # (!always0))))

	.dataa(always0),
	.datab(nRST),
	.datac(always02),
	.datad(\ccif.iwait[0]~1_combout ),
	.cin(gnd),
	.combout(ccifiwait_01),
	.cout());
// synopsys translate_off
defparam \ccif.iwait[0] .lut_mask = 16'hFF4C;
defparam \ccif.iwait[0] .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N24
cycloneive_lcell_comb \ccif.iwait[0]~1 (
// Equation(s):
// \ccif.iwait[0]~1_combout  = ((\nRST~input_o  & ((!always01) # (!LessThan1)))) # (!ccifiwait_0)

	.dataa(LessThan1),
	.datab(ccifiwait_0),
	.datac(nRST),
	.datad(always01),
	.cin(gnd),
	.combout(\ccif.iwait[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ccif.iwait[0]~1 .lut_mask = 16'h73F3;
defparam \ccif.iwait[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
