`include "decode_write_back_if.vh"

module decode_write_back(
	input logic CLK, nRST,
	decode_write_back_if.dw dwif
);

endmodule
