`include "memory_if.vh"

module memory(
	input logic CLK, nRST,
	memory_if.me meif
);

endmodule
