`ifndef COHERENCE_CONTROLLER_IF_VH
`define COHERENCE_CONTROLLER_IF_VH

`include "cpu_types_pkg.vh"
import cpu_types_pkg::*;

interface coherence_controller_if;

	modport cc (
	
	);
endinterface

`endif
